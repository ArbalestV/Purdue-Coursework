module counter
  (
  input wire clk,
  input wire n_reset,
  input wire cnt_up,
  output wire one_k_samples
  );
 /*reg [9:0] data;
 wire clr;*/
 flex_counter #(10) call_counter 
 (.clk(clk),
  .n_rst(n_reset),
  .count_enable(cnt_up),
  .clear(1'b0),//since always cleared up whenever the counter is called
  .rollover_val(10'b1111101000),
  .rollover_flag(one_k_samples)
  );
  //assign clr = one_k_samples;
  
endmodule