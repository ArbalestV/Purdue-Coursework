// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"

// DATE "04/22/2016 22:07:17"

// 
// Device: Altera EP4CE115F29C8 Package FBGA780
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	CLK,
	nRST,
	\syif.halt ,
	\syif.load ,
	\syif.addr ,
	\syif.store ,
	\syif.REN ,
	\syif.WEN ,
	\syif.tbCTRL );
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	CLK;
input 	nRST;
output 	\syif.halt ;
output 	[31:0] \syif.load ;
input 	[31:0] \syif.addr ;
input 	[31:0] \syif.store ;
input 	\syif.REN ;
input 	\syif.WEN ;
input 	\syif.tbCTRL ;

// Design Ports Information
// syif.halt	=>  Location: PIN_AE15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[0]	=>  Location: PIN_T25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[1]	=>  Location: PIN_A17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[2]	=>  Location: PIN_AA15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[3]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[4]	=>  Location: PIN_R27,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[5]	=>  Location: PIN_AB16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[6]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[7]	=>  Location: PIN_J16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[8]	=>  Location: PIN_E17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[9]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[10]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[11]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[12]	=>  Location: PIN_C16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[13]	=>  Location: PIN_G19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[14]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[15]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[16]	=>  Location: PIN_B18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[17]	=>  Location: PIN_H17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[18]	=>  Location: PIN_R23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[19]	=>  Location: PIN_A18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[20]	=>  Location: PIN_Y14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[21]	=>  Location: PIN_AC15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[22]	=>  Location: PIN_J15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[23]	=>  Location: PIN_AD11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[24]	=>  Location: PIN_H16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[25]	=>  Location: PIN_AB14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[26]	=>  Location: PIN_E15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[27]	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[28]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[29]	=>  Location: PIN_AD15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[30]	=>  Location: PIN_G15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[31]	=>  Location: PIN_T21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[1]	=>  Location: PIN_AG15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.tbCTRL	=>  Location: PIN_AH15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[0]	=>  Location: PIN_R24,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[3]	=>  Location: PIN_H13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[2]	=>  Location: PIN_M23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[5]	=>  Location: PIN_A12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[4]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[7]	=>  Location: PIN_F15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[6]	=>  Location: PIN_Y13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[9]	=>  Location: PIN_U3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[8]	=>  Location: PIN_G14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[11]	=>  Location: PIN_A11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[10]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[13]	=>  Location: PIN_D15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[12]	=>  Location: PIN_P26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[15]	=>  Location: PIN_AD14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[14]	=>  Location: PIN_D13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[17]	=>  Location: PIN_AA13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[16]	=>  Location: PIN_B11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[19]	=>  Location: PIN_U4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[18]	=>  Location: PIN_E14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[21]	=>  Location: PIN_D12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[20]	=>  Location: PIN_Y12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[23]	=>  Location: PIN_R7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[22]	=>  Location: PIN_R1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[25]	=>  Location: PIN_F14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[24]	=>  Location: PIN_R2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[27]	=>  Location: PIN_AA12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[26]	=>  Location: PIN_H14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[29]	=>  Location: PIN_C14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[28]	=>  Location: PIN_D14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[31]	=>  Location: PIN_J12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[30]	=>  Location: PIN_C15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.WEN	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.REN	=>  Location: PIN_J14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// nRST	=>  Location: PIN_Y2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// CLK	=>  Location: PIN_J1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[0]	=>  Location: PIN_R26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[1]	=>  Location: PIN_R28,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[2]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[3]	=>  Location: PIN_G21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[4]	=>  Location: PIN_J19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[5]	=>  Location: PIN_H21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[6]	=>  Location: PIN_D16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[7]	=>  Location: PIN_AH18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[8]	=>  Location: PIN_B17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[9]	=>  Location: PIN_AG19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[10]	=>  Location: PIN_P21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[11]	=>  Location: PIN_AH19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[12]	=>  Location: PIN_J17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[13]	=>  Location: PIN_H19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[14]	=>  Location: PIN_R25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[15]	=>  Location: PIN_G18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[16]	=>  Location: PIN_R22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[17]	=>  Location: PIN_T22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[18]	=>  Location: PIN_T26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[19]	=>  Location: PIN_AG18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[20]	=>  Location: PIN_B19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[21]	=>  Location: PIN_Y15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[22]	=>  Location: PIN_G22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[23]	=>  Location: PIN_AB15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[24]	=>  Location: PIN_G20,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[25]	=>  Location: PIN_R21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[26]	=>  Location: PIN_F17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[27]	=>  Location: PIN_J13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[28]	=>  Location: PIN_G16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[29]	=>  Location: PIN_AE17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[30]	=>  Location: PIN_M24,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[31]	=>  Location: PIN_AF17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tms	=>  Location: PIN_P8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tck	=>  Location: PIN_P5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdi	=>  Location: PIN_P7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdo	=>  Location: PIN_P6,	 I/O Standard: 2.5 V,	 Current Strength: Default


wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ;
wire \RAM|LessThan1~0_combout ;
wire \CPU|DP|dWEN_M~q ;
wire \CPU|DP|dREN_M~q ;
wire \ramaddr~0_combout ;
wire \ramaddr~1_combout ;
wire \ramaddr~2_combout ;
wire \ramaddr~3_combout ;
wire \ramaddr~4_combout ;
wire \ramaddr~5_combout ;
wire \ramaddr~6_combout ;
wire \ramaddr~7_combout ;
wire \ramaddr~8_combout ;
wire \ramaddr~9_combout ;
wire \ramaddr~10_combout ;
wire \ramaddr~11_combout ;
wire \ramaddr~12_combout ;
wire \ramaddr~13_combout ;
wire \ramaddr~14_combout ;
wire \ramaddr~15_combout ;
wire \ramaddr~16_combout ;
wire \ramaddr~17_combout ;
wire \ramaddr~18_combout ;
wire \ramaddr~19_combout ;
wire \ramaddr~20_combout ;
wire \ramaddr~21_combout ;
wire \ramaddr~22_combout ;
wire \ramaddr~23_combout ;
wire \ramaddr~24_combout ;
wire \ramaddr~25_combout ;
wire \ramaddr~26_combout ;
wire \ramaddr~27_combout ;
wire \ramaddr~28_combout ;
wire \ramaddr~29_combout ;
wire \ramaddr~30_combout ;
wire \ramaddr~31_combout ;
wire \ramaddr~32_combout ;
wire \ramaddr~33_combout ;
wire \ramaddr~34_combout ;
wire \ramaddr~35_combout ;
wire \ramaddr~36_combout ;
wire \ramaddr~37_combout ;
wire \ramaddr~38_combout ;
wire \ramaddr~39_combout ;
wire \ramaddr~40_combout ;
wire \ramaddr~41_combout ;
wire \ramaddr~42_combout ;
wire \ramaddr~43_combout ;
wire \ramaddr~44_combout ;
wire \ramaddr~45_combout ;
wire \ramaddr~46_combout ;
wire \ramaddr~47_combout ;
wire \ramaddr~48_combout ;
wire \ramaddr~49_combout ;
wire \ramaddr~50_combout ;
wire \ramaddr~51_combout ;
wire \ramaddr~52_combout ;
wire \ramaddr~53_combout ;
wire \ramaddr~54_combout ;
wire \ramaddr~55_combout ;
wire \ramaddr~56_combout ;
wire \ramaddr~57_combout ;
wire \ramaddr~58_combout ;
wire \ramaddr~59_combout ;
wire \ramaddr~60_combout ;
wire \ramaddr~61_combout ;
wire \ramaddr~62_combout ;
wire \ramaddr~63_combout ;
wire \ramWEN~0_combout ;
wire \ramREN~0_combout ;
wire \RAM|always0~21_combout ;
wire \RAM|always1~0_combout ;
wire \RAM|ramif.ramload[0]~0_combout ;
wire \RAM|ramif.ramload[1]~1_combout ;
wire \RAM|ramif.ramload[2]~2_combout ;
wire \RAM|ramif.ramload[3]~3_combout ;
wire \RAM|ramif.ramload[4]~4_combout ;
wire \RAM|ramif.ramload[5]~5_combout ;
wire \RAM|ramif.ramload[6]~6_combout ;
wire \RAM|ramif.ramload[7]~7_combout ;
wire \RAM|ramif.ramload[8]~8_combout ;
wire \RAM|ramif.ramload[9]~9_combout ;
wire \RAM|ramif.ramload[10]~10_combout ;
wire \RAM|ramif.ramload[11]~11_combout ;
wire \RAM|ramif.ramload[12]~12_combout ;
wire \RAM|ramif.ramload[13]~13_combout ;
wire \RAM|ramif.ramload[14]~14_combout ;
wire \RAM|ramif.ramload[15]~15_combout ;
wire \RAM|ramif.ramload[16]~16_combout ;
wire \RAM|ramif.ramload[17]~17_combout ;
wire \RAM|ramif.ramload[18]~18_combout ;
wire \RAM|ramif.ramload[19]~19_combout ;
wire \RAM|ramif.ramload[20]~20_combout ;
wire \RAM|ramif.ramload[21]~21_combout ;
wire \RAM|ramif.ramload[22]~22_combout ;
wire \RAM|ramif.ramload[23]~23_combout ;
wire \RAM|ramif.ramload[24]~24_combout ;
wire \RAM|ramif.ramload[25]~25_combout ;
wire \RAM|ramif.ramload[26]~26_combout ;
wire \RAM|ramif.ramload[27]~27_combout ;
wire \RAM|ramif.ramload[28]~28_combout ;
wire \RAM|ramif.ramload[29]~29_combout ;
wire \RAM|ramif.ramload[30]~30_combout ;
wire \RAM|ramif.ramload[31]~31_combout ;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ;
wire \ramstore~0_combout ;
wire \ramstore~1_combout ;
wire \ramstore~2_combout ;
wire \ramstore~3_combout ;
wire \ramstore~4_combout ;
wire \ramstore~5_combout ;
wire \ramstore~6_combout ;
wire \ramstore~7_combout ;
wire \ramstore~8_combout ;
wire \ramstore~9_combout ;
wire \ramstore~10_combout ;
wire \ramstore~11_combout ;
wire \ramstore~12_combout ;
wire \ramstore~13_combout ;
wire \ramstore~14_combout ;
wire \ramstore~15_combout ;
wire \ramstore~16_combout ;
wire \ramstore~17_combout ;
wire \ramstore~18_combout ;
wire \ramstore~19_combout ;
wire \ramstore~20_combout ;
wire \ramstore~21_combout ;
wire \ramstore~22_combout ;
wire \ramstore~23_combout ;
wire \ramstore~24_combout ;
wire \ramstore~25_combout ;
wire \ramstore~26_combout ;
wire \ramstore~27_combout ;
wire \ramstore~28_combout ;
wire \ramstore~29_combout ;
wire \ramstore~30_combout ;
wire \ramstore~31_combout ;
wire \ramaddr~29_wirecell_combout ;
wire \altera_internal_jtag~TCKUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ;
wire \syif.addr[1]~input_o ;
wire \syif.tbCTRL~input_o ;
wire \syif.addr[0]~input_o ;
wire \syif.addr[3]~input_o ;
wire \syif.addr[2]~input_o ;
wire \syif.addr[5]~input_o ;
wire \syif.addr[4]~input_o ;
wire \syif.addr[7]~input_o ;
wire \syif.addr[6]~input_o ;
wire \syif.addr[9]~input_o ;
wire \syif.addr[8]~input_o ;
wire \syif.addr[11]~input_o ;
wire \syif.addr[10]~input_o ;
wire \syif.addr[13]~input_o ;
wire \syif.addr[12]~input_o ;
wire \syif.addr[15]~input_o ;
wire \syif.addr[14]~input_o ;
wire \syif.addr[17]~input_o ;
wire \syif.addr[16]~input_o ;
wire \syif.addr[19]~input_o ;
wire \syif.addr[18]~input_o ;
wire \syif.addr[21]~input_o ;
wire \syif.addr[20]~input_o ;
wire \syif.addr[23]~input_o ;
wire \syif.addr[22]~input_o ;
wire \syif.addr[25]~input_o ;
wire \syif.addr[24]~input_o ;
wire \syif.addr[27]~input_o ;
wire \syif.addr[26]~input_o ;
wire \syif.addr[29]~input_o ;
wire \syif.addr[28]~input_o ;
wire \syif.addr[31]~input_o ;
wire \syif.addr[30]~input_o ;
wire \syif.WEN~input_o ;
wire \syif.REN~input_o ;
wire \nRST~input_o ;
wire \CLK~input_o ;
wire \syif.store[0]~input_o ;
wire \syif.store[1]~input_o ;
wire \syif.store[2]~input_o ;
wire \syif.store[3]~input_o ;
wire \syif.store[4]~input_o ;
wire \syif.store[5]~input_o ;
wire \syif.store[6]~input_o ;
wire \syif.store[7]~input_o ;
wire \syif.store[8]~input_o ;
wire \syif.store[9]~input_o ;
wire \syif.store[10]~input_o ;
wire \syif.store[11]~input_o ;
wire \syif.store[12]~input_o ;
wire \syif.store[13]~input_o ;
wire \syif.store[14]~input_o ;
wire \syif.store[15]~input_o ;
wire \syif.store[16]~input_o ;
wire \syif.store[17]~input_o ;
wire \syif.store[18]~input_o ;
wire \syif.store[19]~input_o ;
wire \syif.store[20]~input_o ;
wire \syif.store[21]~input_o ;
wire \syif.store[22]~input_o ;
wire \syif.store[23]~input_o ;
wire \syif.store[24]~input_o ;
wire \syif.store[25]~input_o ;
wire \syif.store[26]~input_o ;
wire \syif.store[27]~input_o ;
wire \syif.store[28]~input_o ;
wire \syif.store[29]~input_o ;
wire \syif.store[30]~input_o ;
wire \syif.store[31]~input_o ;
wire \nRST~inputclkctrl_outclk ;
wire \altera_internal_jtag~TCKUTAPclkctrl_outclk ;
wire \CLK~inputclkctrl_outclk ;
wire \CPU|DP|halt_WB~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~10 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg ;
wire [9:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg ;
wire [5:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt ;
wire [15:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR ;
wire [31:0] \CPU|DP|rdata2_M ;
wire [31:0] \CPU|DP|porto_M ;
wire [31:0] \CPU|DP|PROGRAM_COUNTER|pc_out ;
wire [3:0] \RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg ;


ram RAM(
	.is_in_use_reg(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.LessThan1(\RAM|LessThan1~0_combout ),
	.\ramif.ramaddr ({\ramaddr~61_combout ,\ramaddr~63_combout ,\ramaddr~57_combout ,\ramaddr~59_combout ,\ramaddr~53_combout ,\ramaddr~55_combout ,gnd,gnd,gnd,gnd,\ramaddr~41_combout ,\ramaddr~43_combout ,\ramaddr~37_combout ,\ramaddr~39_combout ,\ramaddr~33_combout ,\ramaddr~35_combout ,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\ramaddr~1_combout ,\ramaddr~3_combout }),
	.ramaddr(\ramaddr~5_combout ),
	.ramaddr1(\ramaddr~7_combout ),
	.ramaddr2(\ramaddr~9_combout ),
	.ramaddr3(\ramaddr~11_combout ),
	.ramaddr4(\ramaddr~13_combout ),
	.ramaddr5(\ramaddr~15_combout ),
	.ramaddr6(\ramaddr~17_combout ),
	.ramaddr7(\ramaddr~19_combout ),
	.ramaddr8(\ramaddr~21_combout ),
	.ramaddr9(\ramaddr~23_combout ),
	.ramaddr10(\ramaddr~25_combout ),
	.ramaddr11(\ramaddr~27_combout ),
	.ramaddr12(\ramaddr~29_combout ),
	.ramaddr13(\ramaddr~31_combout ),
	.ramaddr14(\ramaddr~45_combout ),
	.ramaddr15(\ramaddr~47_combout ),
	.ramaddr16(\ramaddr~49_combout ),
	.ramaddr17(\ramaddr~51_combout ),
	.ramWEN(\ramWEN~0_combout ),
	.\ramif.ramREN (\ramREN~0_combout ),
	.always0(\RAM|always0~21_combout ),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~16_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~17_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~18_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~19_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~20_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~21_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~22_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~23_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~24_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~25_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~26_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~27_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~28_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~29_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~30_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~31_combout ),
	.ir_loaded_address_reg_0(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.ir_loaded_address_reg_1(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.ir_loaded_address_reg_2(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.ir_loaded_address_reg_3(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.tdo(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.ramstore(\ramstore~0_combout ),
	.ramstore1(\ramstore~1_combout ),
	.ramstore2(\ramstore~2_combout ),
	.ramstore3(\ramstore~3_combout ),
	.ramstore4(\ramstore~4_combout ),
	.ramstore5(\ramstore~5_combout ),
	.ramstore6(\ramstore~6_combout ),
	.ramstore7(\ramstore~7_combout ),
	.ramstore8(\ramstore~8_combout ),
	.ramstore9(\ramstore~9_combout ),
	.ramstore10(\ramstore~10_combout ),
	.ramstore11(\ramstore~11_combout ),
	.ramstore12(\ramstore~12_combout ),
	.ramstore13(\ramstore~13_combout ),
	.ramstore14(\ramstore~14_combout ),
	.ramstore15(\ramstore~15_combout ),
	.ramstore16(\ramstore~16_combout ),
	.ramstore17(\ramstore~17_combout ),
	.ramstore18(\ramstore~18_combout ),
	.ramstore19(\ramstore~19_combout ),
	.ramstore20(\ramstore~20_combout ),
	.ramstore21(\ramstore~21_combout ),
	.ramstore22(\ramstore~22_combout ),
	.ramstore23(\ramstore~23_combout ),
	.ramstore24(\ramstore~24_combout ),
	.ramstore25(\ramstore~25_combout ),
	.ramstore26(\ramstore~26_combout ),
	.ramstore27(\ramstore~27_combout ),
	.ramstore28(\ramstore~28_combout ),
	.ramstore29(\ramstore~29_combout ),
	.ramstore30(\ramstore~30_combout ),
	.ramstore31(\ramstore~31_combout ),
	.ramaddr18(\ramaddr~29_wirecell_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.irf_reg_0_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.irf_reg_3_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.irf_reg_4_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.node_ena_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.clr_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.virtual_ir_scan_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.state_5(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.state_8(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.nRST(\nRST~input_o ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.altera_internal_jtag1(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.CLK(\CLK~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pipeline CPU(
	.pc_out_3(\CPU|DP|PROGRAM_COUNTER|pc_out [3]),
	.pc_out_2(\CPU|DP|PROGRAM_COUNTER|pc_out [2]),
	.pc_out_5(\CPU|DP|PROGRAM_COUNTER|pc_out [5]),
	.pc_out_4(\CPU|DP|PROGRAM_COUNTER|pc_out [4]),
	.pc_out_7(\CPU|DP|PROGRAM_COUNTER|pc_out [7]),
	.pc_out_6(\CPU|DP|PROGRAM_COUNTER|pc_out [6]),
	.pc_out_9(\CPU|DP|PROGRAM_COUNTER|pc_out [9]),
	.pc_out_8(\CPU|DP|PROGRAM_COUNTER|pc_out [8]),
	.pc_out_11(\CPU|DP|PROGRAM_COUNTER|pc_out [11]),
	.pc_out_10(\CPU|DP|PROGRAM_COUNTER|pc_out [10]),
	.pc_out_13(\CPU|DP|PROGRAM_COUNTER|pc_out [13]),
	.pc_out_12(\CPU|DP|PROGRAM_COUNTER|pc_out [12]),
	.pc_out_15(\CPU|DP|PROGRAM_COUNTER|pc_out [15]),
	.pc_out_14(\CPU|DP|PROGRAM_COUNTER|pc_out [14]),
	.pc_out_17(\CPU|DP|PROGRAM_COUNTER|pc_out [17]),
	.pc_out_16(\CPU|DP|PROGRAM_COUNTER|pc_out [16]),
	.pc_out_19(\CPU|DP|PROGRAM_COUNTER|pc_out [19]),
	.pc_out_18(\CPU|DP|PROGRAM_COUNTER|pc_out [18]),
	.pc_out_21(\CPU|DP|PROGRAM_COUNTER|pc_out [21]),
	.pc_out_20(\CPU|DP|PROGRAM_COUNTER|pc_out [20]),
	.pc_out_23(\CPU|DP|PROGRAM_COUNTER|pc_out [23]),
	.pc_out_22(\CPU|DP|PROGRAM_COUNTER|pc_out [22]),
	.pc_out_25(\CPU|DP|PROGRAM_COUNTER|pc_out [25]),
	.pc_out_24(\CPU|DP|PROGRAM_COUNTER|pc_out [24]),
	.pc_out_27(\CPU|DP|PROGRAM_COUNTER|pc_out [27]),
	.pc_out_26(\CPU|DP|PROGRAM_COUNTER|pc_out [26]),
	.rdata2_M_0(\CPU|DP|rdata2_M [0]),
	.rdata2_M_1(\CPU|DP|rdata2_M [1]),
	.rdata2_M_2(\CPU|DP|rdata2_M [2]),
	.rdata2_M_3(\CPU|DP|rdata2_M [3]),
	.rdata2_M_4(\CPU|DP|rdata2_M [4]),
	.rdata2_M_5(\CPU|DP|rdata2_M [5]),
	.rdata2_M_6(\CPU|DP|rdata2_M [6]),
	.rdata2_M_7(\CPU|DP|rdata2_M [7]),
	.rdata2_M_8(\CPU|DP|rdata2_M [8]),
	.rdata2_M_9(\CPU|DP|rdata2_M [9]),
	.rdata2_M_10(\CPU|DP|rdata2_M [10]),
	.rdata2_M_11(\CPU|DP|rdata2_M [11]),
	.rdata2_M_12(\CPU|DP|rdata2_M [12]),
	.rdata2_M_13(\CPU|DP|rdata2_M [13]),
	.rdata2_M_14(\CPU|DP|rdata2_M [14]),
	.rdata2_M_15(\CPU|DP|rdata2_M [15]),
	.rdata2_M_16(\CPU|DP|rdata2_M [16]),
	.rdata2_M_17(\CPU|DP|rdata2_M [17]),
	.rdata2_M_18(\CPU|DP|rdata2_M [18]),
	.rdata2_M_19(\CPU|DP|rdata2_M [19]),
	.rdata2_M_20(\CPU|DP|rdata2_M [20]),
	.rdata2_M_21(\CPU|DP|rdata2_M [21]),
	.rdata2_M_22(\CPU|DP|rdata2_M [22]),
	.rdata2_M_23(\CPU|DP|rdata2_M [23]),
	.rdata2_M_24(\CPU|DP|rdata2_M [24]),
	.rdata2_M_25(\CPU|DP|rdata2_M [25]),
	.rdata2_M_26(\CPU|DP|rdata2_M [26]),
	.rdata2_M_27(\CPU|DP|rdata2_M [27]),
	.rdata2_M_28(\CPU|DP|rdata2_M [28]),
	.rdata2_M_29(\CPU|DP|rdata2_M [29]),
	.rdata2_M_30(\CPU|DP|rdata2_M [30]),
	.rdata2_M_31(\CPU|DP|rdata2_M [31]),
	.LessThan1(\RAM|LessThan1~0_combout ),
	.porto_M_1(\CPU|DP|porto_M [1]),
	.pc_out_1(\CPU|DP|PROGRAM_COUNTER|pc_out [1]),
	.dWEN_M(\CPU|DP|dWEN_M~q ),
	.dREN_M(\CPU|DP|dREN_M~q ),
	.porto_M_0(\CPU|DP|porto_M [0]),
	.pc_out_0(\CPU|DP|PROGRAM_COUNTER|pc_out [0]),
	.porto_M_3(\CPU|DP|porto_M [3]),
	.porto_M_2(\CPU|DP|porto_M [2]),
	.porto_M_5(\CPU|DP|porto_M [5]),
	.porto_M_4(\CPU|DP|porto_M [4]),
	.porto_M_7(\CPU|DP|porto_M [7]),
	.porto_M_6(\CPU|DP|porto_M [6]),
	.porto_M_9(\CPU|DP|porto_M [9]),
	.porto_M_8(\CPU|DP|porto_M [8]),
	.porto_M_11(\CPU|DP|porto_M [11]),
	.porto_M_10(\CPU|DP|porto_M [10]),
	.porto_M_13(\CPU|DP|porto_M [13]),
	.porto_M_12(\CPU|DP|porto_M [12]),
	.porto_M_15(\CPU|DP|porto_M [15]),
	.porto_M_14(\CPU|DP|porto_M [14]),
	.porto_M_17(\CPU|DP|porto_M [17]),
	.porto_M_16(\CPU|DP|porto_M [16]),
	.porto_M_19(\CPU|DP|porto_M [19]),
	.porto_M_18(\CPU|DP|porto_M [18]),
	.porto_M_21(\CPU|DP|porto_M [21]),
	.porto_M_20(\CPU|DP|porto_M [20]),
	.porto_M_23(\CPU|DP|porto_M [23]),
	.porto_M_22(\CPU|DP|porto_M [22]),
	.porto_M_25(\CPU|DP|porto_M [25]),
	.porto_M_24(\CPU|DP|porto_M [24]),
	.porto_M_27(\CPU|DP|porto_M [27]),
	.porto_M_26(\CPU|DP|porto_M [26]),
	.porto_M_29(\CPU|DP|porto_M [29]),
	.pc_out_29(\CPU|DP|PROGRAM_COUNTER|pc_out [29]),
	.porto_M_28(\CPU|DP|porto_M [28]),
	.pc_out_28(\CPU|DP|PROGRAM_COUNTER|pc_out [28]),
	.porto_M_31(\CPU|DP|porto_M [31]),
	.pc_out_31(\CPU|DP|PROGRAM_COUNTER|pc_out [31]),
	.porto_M_30(\CPU|DP|porto_M [30]),
	.pc_out_30(\CPU|DP|PROGRAM_COUNTER|pc_out [30]),
	.always0(\RAM|always0~21_combout ),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~16_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~17_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~18_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~19_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~20_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~21_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~22_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~23_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~24_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~25_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~26_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~27_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~28_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~29_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~30_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~31_combout ),
	.nRST(\nRST~input_o ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.CLK(\CLK~inputclkctrl_outclk ),
	.halt_WB(\CPU|DP|halt_WB~q ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X53_Y35_N12
cycloneive_lcell_comb \ramaddr~0 (
// Equation(s):
// \ramaddr~0_combout  = (dWEN_M1 & (porto_M_1)) # (!dWEN_M1 & ((dREN_M1 & (porto_M_1)) # (!dREN_M1 & ((pc_out_1)))))

	.dataa(\CPU|DP|dWEN_M~q ),
	.datab(\CPU|DP|porto_M [1]),
	.datac(\CPU|DP|PROGRAM_COUNTER|pc_out [1]),
	.datad(\CPU|DP|dREN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~0 .lut_mask = 16'hCCD8;
defparam \ramaddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N30
cycloneive_lcell_comb \ramaddr~1 (
// Equation(s):
// \ramaddr~1_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[1]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~0_combout )))

	.dataa(gnd),
	.datab(\syif.addr[1]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~0_combout ),
	.cin(gnd),
	.combout(\ramaddr~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~1 .lut_mask = 16'hCFC0;
defparam \ramaddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N16
cycloneive_lcell_comb \ramaddr~2 (
// Equation(s):
// \ramaddr~2_combout  = (dREN_M1 & (((porto_M_0)))) # (!dREN_M1 & ((dWEN_M1 & ((porto_M_0))) # (!dWEN_M1 & (pc_out_0))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [0]),
	.datab(\CPU|DP|dREN_M~q ),
	.datac(\CPU|DP|dWEN_M~q ),
	.datad(\CPU|DP|porto_M [0]),
	.cin(gnd),
	.combout(\ramaddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~2 .lut_mask = 16'hFE02;
defparam \ramaddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N20
cycloneive_lcell_comb \ramaddr~3 (
// Equation(s):
// \ramaddr~3_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~2_combout )))

	.dataa(gnd),
	.datab(\syif.addr[0]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~2_combout ),
	.cin(gnd),
	.combout(\ramaddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~3 .lut_mask = 16'hCFC0;
defparam \ramaddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N16
cycloneive_lcell_comb \ramaddr~4 (
// Equation(s):
// \ramaddr~4_combout  = (dREN_M1 & (((porto_M_3)))) # (!dREN_M1 & ((dWEN_M1 & (porto_M_3)) # (!dWEN_M1 & ((pc_out_3)))))

	.dataa(\CPU|DP|dREN_M~q ),
	.datab(\CPU|DP|dWEN_M~q ),
	.datac(\CPU|DP|porto_M [3]),
	.datad(\CPU|DP|PROGRAM_COUNTER|pc_out [3]),
	.cin(gnd),
	.combout(\ramaddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~4 .lut_mask = 16'hF1E0;
defparam \ramaddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N0
cycloneive_lcell_comb \ramaddr~5 (
// Equation(s):
// \ramaddr~5_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[3]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~4_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[3]~input_o ),
	.datac(\ramaddr~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~5 .lut_mask = 16'hD8D8;
defparam \ramaddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N2
cycloneive_lcell_comb \ramaddr~6 (
// Equation(s):
// \ramaddr~6_combout  = (dREN_M1 & (porto_M_2)) # (!dREN_M1 & ((dWEN_M1 & (porto_M_2)) # (!dWEN_M1 & ((pc_out_2)))))

	.dataa(\CPU|DP|dREN_M~q ),
	.datab(\CPU|DP|porto_M [2]),
	.datac(\CPU|DP|dWEN_M~q ),
	.datad(\CPU|DP|PROGRAM_COUNTER|pc_out [2]),
	.cin(gnd),
	.combout(\ramaddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~6 .lut_mask = 16'hCDC8;
defparam \ramaddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N2
cycloneive_lcell_comb \ramaddr~7 (
// Equation(s):
// \ramaddr~7_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[2]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~6_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[2]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~6_combout ),
	.cin(gnd),
	.combout(\ramaddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~7 .lut_mask = 16'hDD88;
defparam \ramaddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N14
cycloneive_lcell_comb \ramaddr~8 (
// Equation(s):
// \ramaddr~8_combout  = (dREN_M1 & (((porto_M_5)))) # (!dREN_M1 & ((dWEN_M1 & ((porto_M_5))) # (!dWEN_M1 & (pc_out_5))))

	.dataa(\CPU|DP|dREN_M~q ),
	.datab(\CPU|DP|PROGRAM_COUNTER|pc_out [5]),
	.datac(\CPU|DP|porto_M [5]),
	.datad(\CPU|DP|dWEN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~8 .lut_mask = 16'hF0E4;
defparam \ramaddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N22
cycloneive_lcell_comb \ramaddr~9 (
// Equation(s):
// \ramaddr~9_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~8_combout )))

	.dataa(gnd),
	.datab(\syif.addr[5]~input_o ),
	.datac(\ramaddr~8_combout ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~9 .lut_mask = 16'hCCF0;
defparam \ramaddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N28
cycloneive_lcell_comb \ramaddr~10 (
// Equation(s):
// \ramaddr~10_combout  = (dWEN_M1 & (porto_M_4)) # (!dWEN_M1 & ((dREN_M1 & (porto_M_4)) # (!dREN_M1 & ((pc_out_4)))))

	.dataa(\CPU|DP|dWEN_M~q ),
	.datab(\CPU|DP|porto_M [4]),
	.datac(\CPU|DP|dREN_M~q ),
	.datad(\CPU|DP|PROGRAM_COUNTER|pc_out [4]),
	.cin(gnd),
	.combout(\ramaddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~10 .lut_mask = 16'hCDC8;
defparam \ramaddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N16
cycloneive_lcell_comb \ramaddr~11 (
// Equation(s):
// \ramaddr~11_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[4]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~10_combout )))

	.dataa(\syif.addr[4]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~10_combout ),
	.cin(gnd),
	.combout(\ramaddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~11 .lut_mask = 16'hBB88;
defparam \ramaddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N10
cycloneive_lcell_comb \ramaddr~12 (
// Equation(s):
// \ramaddr~12_combout  = (dWEN_M1 & (((porto_M_7)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_7))) # (!dREN_M1 & (pc_out_7))))

	.dataa(\CPU|DP|dWEN_M~q ),
	.datab(\CPU|DP|PROGRAM_COUNTER|pc_out [7]),
	.datac(\CPU|DP|porto_M [7]),
	.datad(\CPU|DP|dREN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~12 .lut_mask = 16'hF0E4;
defparam \ramaddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N26
cycloneive_lcell_comb \ramaddr~13 (
// Equation(s):
// \ramaddr~13_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~12_combout )))

	.dataa(gnd),
	.datab(\syif.addr[7]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~12_combout ),
	.cin(gnd),
	.combout(\ramaddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~13 .lut_mask = 16'hCFC0;
defparam \ramaddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N18
cycloneive_lcell_comb \ramaddr~14 (
// Equation(s):
// \ramaddr~14_combout  = (dWEN_M1 & (((porto_M_6)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_6))) # (!dREN_M1 & (pc_out_6))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [6]),
	.datab(\CPU|DP|dWEN_M~q ),
	.datac(\CPU|DP|dREN_M~q ),
	.datad(\CPU|DP|porto_M [6]),
	.cin(gnd),
	.combout(\ramaddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~14 .lut_mask = 16'hFE02;
defparam \ramaddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N28
cycloneive_lcell_comb \ramaddr~15 (
// Equation(s):
// \ramaddr~15_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[6]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~14_combout )))

	.dataa(gnd),
	.datab(\syif.addr[6]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~14_combout ),
	.cin(gnd),
	.combout(\ramaddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~15 .lut_mask = 16'hCFC0;
defparam \ramaddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N28
cycloneive_lcell_comb \ramaddr~16 (
// Equation(s):
// \ramaddr~16_combout  = (dWEN_M1 & (((porto_M_9)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_9))) # (!dREN_M1 & (pc_out_9))))

	.dataa(\CPU|DP|dWEN_M~q ),
	.datab(\CPU|DP|PROGRAM_COUNTER|pc_out [9]),
	.datac(\CPU|DP|porto_M [9]),
	.datad(\CPU|DP|dREN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~16 .lut_mask = 16'hF0E4;
defparam \ramaddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N26
cycloneive_lcell_comb \ramaddr~17 (
// Equation(s):
// \ramaddr~17_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[9]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~16_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[9]~input_o ),
	.datad(\ramaddr~16_combout ),
	.cin(gnd),
	.combout(\ramaddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~17 .lut_mask = 16'hF3C0;
defparam \ramaddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N16
cycloneive_lcell_comb \ramaddr~18 (
// Equation(s):
// \ramaddr~18_combout  = (dREN_M1 & (((porto_M_8)))) # (!dREN_M1 & ((dWEN_M1 & ((porto_M_8))) # (!dWEN_M1 & (pc_out_8))))

	.dataa(\CPU|DP|dREN_M~q ),
	.datab(\CPU|DP|PROGRAM_COUNTER|pc_out [8]),
	.datac(\CPU|DP|dWEN_M~q ),
	.datad(\CPU|DP|porto_M [8]),
	.cin(gnd),
	.combout(\ramaddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~18 .lut_mask = 16'hFE04;
defparam \ramaddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N20
cycloneive_lcell_comb \ramaddr~19 (
// Equation(s):
// \ramaddr~19_combout  = (\syif.tbCTRL~input_o  & ((\syif.addr[8]~input_o ))) # (!\syif.tbCTRL~input_o  & (\ramaddr~18_combout ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~18_combout ),
	.datad(\syif.addr[8]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~19 .lut_mask = 16'hFC30;
defparam \ramaddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N22
cycloneive_lcell_comb \ramaddr~20 (
// Equation(s):
// \ramaddr~20_combout  = (dWEN_M1 & (((porto_M_11)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_11))) # (!dREN_M1 & (pc_out_11))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [11]),
	.datab(\CPU|DP|dWEN_M~q ),
	.datac(\CPU|DP|porto_M [11]),
	.datad(\CPU|DP|dREN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~20 .lut_mask = 16'hF0E2;
defparam \ramaddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N18
cycloneive_lcell_comb \ramaddr~21 (
// Equation(s):
// \ramaddr~21_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~20_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[11]~input_o ),
	.datad(\ramaddr~20_combout ),
	.cin(gnd),
	.combout(\ramaddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~21 .lut_mask = 16'hF5A0;
defparam \ramaddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N18
cycloneive_lcell_comb \ramaddr~22 (
// Equation(s):
// \ramaddr~22_combout  = (dWEN_M1 & (porto_M_10)) # (!dWEN_M1 & ((dREN_M1 & (porto_M_10)) # (!dREN_M1 & ((pc_out_10)))))

	.dataa(\CPU|DP|dWEN_M~q ),
	.datab(\CPU|DP|porto_M [10]),
	.datac(\CPU|DP|PROGRAM_COUNTER|pc_out [10]),
	.datad(\CPU|DP|dREN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~22 .lut_mask = 16'hCCD8;
defparam \ramaddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N24
cycloneive_lcell_comb \ramaddr~23 (
// Equation(s):
// \ramaddr~23_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~22_combout )))

	.dataa(\syif.addr[10]~input_o ),
	.datab(\ramaddr~22_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~23 .lut_mask = 16'hACAC;
defparam \ramaddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N14
cycloneive_lcell_comb \ramaddr~24 (
// Equation(s):
// \ramaddr~24_combout  = (dWEN_M1 & (((porto_M_13)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_13))) # (!dREN_M1 & (pc_out_13))))

	.dataa(\CPU|DP|dWEN_M~q ),
	.datab(\CPU|DP|dREN_M~q ),
	.datac(\CPU|DP|PROGRAM_COUNTER|pc_out [13]),
	.datad(\CPU|DP|porto_M [13]),
	.cin(gnd),
	.combout(\ramaddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~24 .lut_mask = 16'hFE10;
defparam \ramaddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N16
cycloneive_lcell_comb \ramaddr~25 (
// Equation(s):
// \ramaddr~25_combout  = (\syif.tbCTRL~input_o  & ((\syif.addr[13]~input_o ))) # (!\syif.tbCTRL~input_o  & (\ramaddr~24_combout ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\ramaddr~24_combout ),
	.datad(\syif.addr[13]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~25 .lut_mask = 16'hFA50;
defparam \ramaddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N24
cycloneive_lcell_comb \ramaddr~26 (
// Equation(s):
// \ramaddr~26_combout  = (dREN_M1 & (((porto_M_12)))) # (!dREN_M1 & ((dWEN_M1 & ((porto_M_12))) # (!dWEN_M1 & (pc_out_12))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [12]),
	.datab(\CPU|DP|dREN_M~q ),
	.datac(\CPU|DP|dWEN_M~q ),
	.datad(\CPU|DP|porto_M [12]),
	.cin(gnd),
	.combout(\ramaddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~26 .lut_mask = 16'hFE02;
defparam \ramaddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N28
cycloneive_lcell_comb \ramaddr~27 (
// Equation(s):
// \ramaddr~27_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[12]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~26_combout )))

	.dataa(\syif.addr[12]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~26_combout ),
	.cin(gnd),
	.combout(\ramaddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~27 .lut_mask = 16'hAFA0;
defparam \ramaddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N2
cycloneive_lcell_comb \ramaddr~28 (
// Equation(s):
// \ramaddr~28_combout  = (dREN_M1 & (((porto_M_15)))) # (!dREN_M1 & ((dWEN_M1 & ((porto_M_15))) # (!dWEN_M1 & (pc_out_15))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [15]),
	.datab(\CPU|DP|dREN_M~q ),
	.datac(\CPU|DP|dWEN_M~q ),
	.datad(\CPU|DP|porto_M [15]),
	.cin(gnd),
	.combout(\ramaddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~28 .lut_mask = 16'hFE02;
defparam \ramaddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N4
cycloneive_lcell_comb \ramaddr~29 (
// Equation(s):
// \ramaddr~29_combout  = (\syif.tbCTRL~input_o  & (!\syif.addr[15]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~28_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[15]~input_o ),
	.datad(\ramaddr~28_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29 .lut_mask = 16'h0C3F;
defparam \ramaddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N20
cycloneive_lcell_comb \ramaddr~30 (
// Equation(s):
// \ramaddr~30_combout  = (dREN_M1 & (((porto_M_14)))) # (!dREN_M1 & ((dWEN_M1 & (porto_M_14)) # (!dWEN_M1 & ((pc_out_14)))))

	.dataa(\CPU|DP|dREN_M~q ),
	.datab(\CPU|DP|dWEN_M~q ),
	.datac(\CPU|DP|porto_M [14]),
	.datad(\CPU|DP|PROGRAM_COUNTER|pc_out [14]),
	.cin(gnd),
	.combout(\ramaddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~30 .lut_mask = 16'hF1E0;
defparam \ramaddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N28
cycloneive_lcell_comb \ramaddr~31 (
// Equation(s):
// \ramaddr~31_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~30_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[14]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~30_combout ),
	.cin(gnd),
	.combout(\ramaddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~31 .lut_mask = 16'hDD88;
defparam \ramaddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N28
cycloneive_lcell_comb \ramaddr~32 (
// Equation(s):
// \ramaddr~32_combout  = (dWEN_M1 & (porto_M_17)) # (!dWEN_M1 & ((dREN_M1 & (porto_M_17)) # (!dREN_M1 & ((pc_out_17)))))

	.dataa(\CPU|DP|porto_M [17]),
	.datab(\CPU|DP|dWEN_M~q ),
	.datac(\CPU|DP|dREN_M~q ),
	.datad(\CPU|DP|PROGRAM_COUNTER|pc_out [17]),
	.cin(gnd),
	.combout(\ramaddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~32 .lut_mask = 16'hABA8;
defparam \ramaddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N24
cycloneive_lcell_comb \ramaddr~33 (
// Equation(s):
// \ramaddr~33_combout  = (\syif.tbCTRL~input_o  & ((\syif.addr[17]~input_o ))) # (!\syif.tbCTRL~input_o  & (\ramaddr~32_combout ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~32_combout ),
	.datad(\syif.addr[17]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~33 .lut_mask = 16'hFC30;
defparam \ramaddr~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N6
cycloneive_lcell_comb \ramaddr~34 (
// Equation(s):
// \ramaddr~34_combout  = (dREN_M1 & (porto_M_16)) # (!dREN_M1 & ((dWEN_M1 & (porto_M_16)) # (!dWEN_M1 & ((pc_out_16)))))

	.dataa(\CPU|DP|dREN_M~q ),
	.datab(\CPU|DP|porto_M [16]),
	.datac(\CPU|DP|PROGRAM_COUNTER|pc_out [16]),
	.datad(\CPU|DP|dWEN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~34 .lut_mask = 16'hCCD8;
defparam \ramaddr~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N10
cycloneive_lcell_comb \ramaddr~35 (
// Equation(s):
// \ramaddr~35_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[16]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~34_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[16]~input_o ),
	.datad(\ramaddr~34_combout ),
	.cin(gnd),
	.combout(\ramaddr~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~35 .lut_mask = 16'hF3C0;
defparam \ramaddr~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N24
cycloneive_lcell_comb \ramaddr~36 (
// Equation(s):
// \ramaddr~36_combout  = (dWEN_M1 & (((porto_M_19)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_19))) # (!dREN_M1 & (pc_out_19))))

	.dataa(\CPU|DP|dWEN_M~q ),
	.datab(\CPU|DP|dREN_M~q ),
	.datac(\CPU|DP|PROGRAM_COUNTER|pc_out [19]),
	.datad(\CPU|DP|porto_M [19]),
	.cin(gnd),
	.combout(\ramaddr~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~36 .lut_mask = 16'hFE10;
defparam \ramaddr~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N2
cycloneive_lcell_comb \ramaddr~37 (
// Equation(s):
// \ramaddr~37_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~36_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[19]~input_o ),
	.datad(\ramaddr~36_combout ),
	.cin(gnd),
	.combout(\ramaddr~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~37 .lut_mask = 16'hF5A0;
defparam \ramaddr~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N4
cycloneive_lcell_comb \ramaddr~38 (
// Equation(s):
// \ramaddr~38_combout  = (dREN_M1 & (((porto_M_18)))) # (!dREN_M1 & ((dWEN_M1 & ((porto_M_18))) # (!dWEN_M1 & (pc_out_18))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [18]),
	.datab(\CPU|DP|porto_M [18]),
	.datac(\CPU|DP|dREN_M~q ),
	.datad(\CPU|DP|dWEN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~38 .lut_mask = 16'hCCCA;
defparam \ramaddr~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N4
cycloneive_lcell_comb \ramaddr~39 (
// Equation(s):
// \ramaddr~39_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~38_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[18]~input_o ),
	.datad(\ramaddr~38_combout ),
	.cin(gnd),
	.combout(\ramaddr~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~39 .lut_mask = 16'hF5A0;
defparam \ramaddr~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N14
cycloneive_lcell_comb \ramaddr~40 (
// Equation(s):
// \ramaddr~40_combout  = (dWEN_M1 & (((porto_M_21)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_21))) # (!dREN_M1 & (pc_out_21))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [21]),
	.datab(\CPU|DP|dWEN_M~q ),
	.datac(\CPU|DP|dREN_M~q ),
	.datad(\CPU|DP|porto_M [21]),
	.cin(gnd),
	.combout(\ramaddr~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~40 .lut_mask = 16'hFE02;
defparam \ramaddr~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N4
cycloneive_lcell_comb \ramaddr~41 (
// Equation(s):
// \ramaddr~41_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[21]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~40_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[21]~input_o ),
	.datad(\ramaddr~40_combout ),
	.cin(gnd),
	.combout(\ramaddr~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~41 .lut_mask = 16'hF3C0;
defparam \ramaddr~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N18
cycloneive_lcell_comb \ramaddr~42 (
// Equation(s):
// \ramaddr~42_combout  = (dREN_M1 & (((porto_M_20)))) # (!dREN_M1 & ((dWEN_M1 & ((porto_M_20))) # (!dWEN_M1 & (pc_out_20))))

	.dataa(\CPU|DP|dREN_M~q ),
	.datab(\CPU|DP|PROGRAM_COUNTER|pc_out [20]),
	.datac(\CPU|DP|porto_M [20]),
	.datad(\CPU|DP|dWEN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~42 .lut_mask = 16'hF0E4;
defparam \ramaddr~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N2
cycloneive_lcell_comb \ramaddr~43 (
// Equation(s):
// \ramaddr~43_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~42_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[20]~input_o ),
	.datad(\ramaddr~42_combout ),
	.cin(gnd),
	.combout(\ramaddr~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~43 .lut_mask = 16'hF3C0;
defparam \ramaddr~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N2
cycloneive_lcell_comb \ramaddr~44 (
// Equation(s):
// \ramaddr~44_combout  = (dWEN_M1 & (((porto_M_23)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_23))) # (!dREN_M1 & (pc_out_23))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [23]),
	.datab(\CPU|DP|porto_M [23]),
	.datac(\CPU|DP|dWEN_M~q ),
	.datad(\CPU|DP|dREN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~44 .lut_mask = 16'hCCCA;
defparam \ramaddr~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N4
cycloneive_lcell_comb \ramaddr~45 (
// Equation(s):
// \ramaddr~45_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[23]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~44_combout )))

	.dataa(gnd),
	.datab(\syif.addr[23]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~44_combout ),
	.cin(gnd),
	.combout(\ramaddr~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~45 .lut_mask = 16'hCFC0;
defparam \ramaddr~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N20
cycloneive_lcell_comb \ramaddr~46 (
// Equation(s):
// \ramaddr~46_combout  = (dWEN_M1 & (((porto_M_22)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_22))) # (!dREN_M1 & (pc_out_22))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [22]),
	.datab(\CPU|DP|porto_M [22]),
	.datac(\CPU|DP|dWEN_M~q ),
	.datad(\CPU|DP|dREN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~46 .lut_mask = 16'hCCCA;
defparam \ramaddr~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N2
cycloneive_lcell_comb \ramaddr~47 (
// Equation(s):
// \ramaddr~47_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[22]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~46_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[22]~input_o ),
	.datac(\ramaddr~46_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~47 .lut_mask = 16'hD8D8;
defparam \ramaddr~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N22
cycloneive_lcell_comb \ramaddr~48 (
// Equation(s):
// \ramaddr~48_combout  = (dREN_M1 & (porto_M_25)) # (!dREN_M1 & ((dWEN_M1 & (porto_M_25)) # (!dWEN_M1 & ((pc_out_25)))))

	.dataa(\CPU|DP|dREN_M~q ),
	.datab(\CPU|DP|porto_M [25]),
	.datac(\CPU|DP|dWEN_M~q ),
	.datad(\CPU|DP|PROGRAM_COUNTER|pc_out [25]),
	.cin(gnd),
	.combout(\ramaddr~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~48 .lut_mask = 16'hCDC8;
defparam \ramaddr~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N28
cycloneive_lcell_comb \ramaddr~49 (
// Equation(s):
// \ramaddr~49_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[25]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~48_combout )))

	.dataa(gnd),
	.datab(\syif.addr[25]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~48_combout ),
	.cin(gnd),
	.combout(\ramaddr~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~49 .lut_mask = 16'hCFC0;
defparam \ramaddr~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N10
cycloneive_lcell_comb \ramaddr~50 (
// Equation(s):
// \ramaddr~50_combout  = (dWEN_M1 & (((porto_M_24)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_24))) # (!dREN_M1 & (pc_out_24))))

	.dataa(\CPU|DP|dWEN_M~q ),
	.datab(\CPU|DP|dREN_M~q ),
	.datac(\CPU|DP|PROGRAM_COUNTER|pc_out [24]),
	.datad(\CPU|DP|porto_M [24]),
	.cin(gnd),
	.combout(\ramaddr~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~50 .lut_mask = 16'hFE10;
defparam \ramaddr~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N8
cycloneive_lcell_comb \ramaddr~51 (
// Equation(s):
// \ramaddr~51_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~50_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[24]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~50_combout ),
	.cin(gnd),
	.combout(\ramaddr~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~51 .lut_mask = 16'hDD88;
defparam \ramaddr~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N2
cycloneive_lcell_comb \ramaddr~52 (
// Equation(s):
// \ramaddr~52_combout  = (dWEN_M1 & (porto_M_27)) # (!dWEN_M1 & ((dREN_M1 & (porto_M_27)) # (!dREN_M1 & ((pc_out_27)))))

	.dataa(\CPU|DP|porto_M [27]),
	.datab(\CPU|DP|dWEN_M~q ),
	.datac(\CPU|DP|dREN_M~q ),
	.datad(\CPU|DP|PROGRAM_COUNTER|pc_out [27]),
	.cin(gnd),
	.combout(\ramaddr~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~52 .lut_mask = 16'hABA8;
defparam \ramaddr~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N8
cycloneive_lcell_comb \ramaddr~53 (
// Equation(s):
// \ramaddr~53_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~52_combout )))

	.dataa(\syif.addr[27]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~52_combout ),
	.cin(gnd),
	.combout(\ramaddr~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~53 .lut_mask = 16'hAFA0;
defparam \ramaddr~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N16
cycloneive_lcell_comb \ramaddr~54 (
// Equation(s):
// \ramaddr~54_combout  = (dREN_M1 & (((porto_M_26)))) # (!dREN_M1 & ((dWEN_M1 & ((porto_M_26))) # (!dWEN_M1 & (pc_out_26))))

	.dataa(\CPU|DP|dREN_M~q ),
	.datab(\CPU|DP|PROGRAM_COUNTER|pc_out [26]),
	.datac(\CPU|DP|porto_M [26]),
	.datad(\CPU|DP|dWEN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~54 .lut_mask = 16'hF0E4;
defparam \ramaddr~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N30
cycloneive_lcell_comb \ramaddr~55 (
// Equation(s):
// \ramaddr~55_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~54_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[26]~input_o ),
	.datad(\ramaddr~54_combout ),
	.cin(gnd),
	.combout(\ramaddr~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~55 .lut_mask = 16'hF3C0;
defparam \ramaddr~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N6
cycloneive_lcell_comb \ramaddr~56 (
// Equation(s):
// \ramaddr~56_combout  = (dWEN_M1 & (((porto_M_29)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_29))) # (!dREN_M1 & (pc_out_29))))

	.dataa(\CPU|DP|dWEN_M~q ),
	.datab(\CPU|DP|PROGRAM_COUNTER|pc_out [29]),
	.datac(\CPU|DP|dREN_M~q ),
	.datad(\CPU|DP|porto_M [29]),
	.cin(gnd),
	.combout(\ramaddr~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~56 .lut_mask = 16'hFE04;
defparam \ramaddr~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N24
cycloneive_lcell_comb \ramaddr~57 (
// Equation(s):
// \ramaddr~57_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[29]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~56_combout )))

	.dataa(\syif.addr[29]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~56_combout ),
	.cin(gnd),
	.combout(\ramaddr~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~57 .lut_mask = 16'hBB88;
defparam \ramaddr~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N12
cycloneive_lcell_comb \ramaddr~58 (
// Equation(s):
// \ramaddr~58_combout  = (dWEN_M1 & (((porto_M_28)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_28))) # (!dREN_M1 & (pc_out_28))))

	.dataa(\CPU|DP|dWEN_M~q ),
	.datab(\CPU|DP|PROGRAM_COUNTER|pc_out [28]),
	.datac(\CPU|DP|dREN_M~q ),
	.datad(\CPU|DP|porto_M [28]),
	.cin(gnd),
	.combout(\ramaddr~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~58 .lut_mask = 16'hFE04;
defparam \ramaddr~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N14
cycloneive_lcell_comb \ramaddr~59 (
// Equation(s):
// \ramaddr~59_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~58_combout )))

	.dataa(gnd),
	.datab(\syif.addr[28]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~58_combout ),
	.cin(gnd),
	.combout(\ramaddr~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~59 .lut_mask = 16'hCFC0;
defparam \ramaddr~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N6
cycloneive_lcell_comb \ramaddr~60 (
// Equation(s):
// \ramaddr~60_combout  = (dREN_M1 & (((porto_M_31)))) # (!dREN_M1 & ((dWEN_M1 & ((porto_M_31))) # (!dWEN_M1 & (pc_out_31))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [31]),
	.datab(\CPU|DP|dREN_M~q ),
	.datac(\CPU|DP|dWEN_M~q ),
	.datad(\CPU|DP|porto_M [31]),
	.cin(gnd),
	.combout(\ramaddr~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~60 .lut_mask = 16'hFE02;
defparam \ramaddr~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N8
cycloneive_lcell_comb \ramaddr~61 (
// Equation(s):
// \ramaddr~61_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~60_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[31]~input_o ),
	.datad(\ramaddr~60_combout ),
	.cin(gnd),
	.combout(\ramaddr~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~61 .lut_mask = 16'hF3C0;
defparam \ramaddr~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N24
cycloneive_lcell_comb \ramaddr~62 (
// Equation(s):
// \ramaddr~62_combout  = (dWEN_M1 & (((porto_M_30)))) # (!dWEN_M1 & ((dREN_M1 & ((porto_M_30))) # (!dREN_M1 & (pc_out_30))))

	.dataa(\CPU|DP|PROGRAM_COUNTER|pc_out [30]),
	.datab(\CPU|DP|dWEN_M~q ),
	.datac(\CPU|DP|porto_M [30]),
	.datad(\CPU|DP|dREN_M~q ),
	.cin(gnd),
	.combout(\ramaddr~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~62 .lut_mask = 16'hF0E2;
defparam \ramaddr~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N18
cycloneive_lcell_comb \ramaddr~63 (
// Equation(s):
// \ramaddr~63_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[30]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~62_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[30]~input_o ),
	.datad(\ramaddr~62_combout ),
	.cin(gnd),
	.combout(\ramaddr~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~63 .lut_mask = 16'hF3C0;
defparam \ramaddr~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N22
cycloneive_lcell_comb \ramWEN~0 (
// Equation(s):
// \ramWEN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.WEN~input_o )) # (!\syif.tbCTRL~input_o  & ((!dWEN_M1)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.WEN~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|dWEN_M~q ),
	.cin(gnd),
	.combout(\ramWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramWEN~0 .lut_mask = 16'h2277;
defparam \ramWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N12
cycloneive_lcell_comb \ramREN~0 (
// Equation(s):
// \ramREN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.REN~input_o )) # (!\syif.tbCTRL~input_o  & ((dWEN_M1)))

	.dataa(gnd),
	.datab(\syif.REN~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|dWEN_M~q ),
	.cin(gnd),
	.combout(\ramREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~0 .lut_mask = 16'h3F30;
defparam \ramREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N14
cycloneive_lcell_comb \ramstore~0 (
// Equation(s):
// \ramstore~0_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[0]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_0))

	.dataa(\CPU|DP|rdata2_M [0]),
	.datab(\syif.store[0]~input_o ),
	.datac(gnd),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~0 .lut_mask = 16'hCCAA;
defparam \ramstore~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N0
cycloneive_lcell_comb \ramstore~1 (
// Equation(s):
// \ramstore~1_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[1]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_1))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rdata2_M [1]),
	.datad(\syif.store[1]~input_o ),
	.cin(gnd),
	.combout(\ramstore~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~1 .lut_mask = 16'hFC30;
defparam \ramstore~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N22
cycloneive_lcell_comb \ramstore~2 (
// Equation(s):
// \ramstore~2_combout  = (\syif.tbCTRL~input_o  & (\syif.store[2]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_2)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[2]~input_o ),
	.datad(\CPU|DP|rdata2_M [2]),
	.cin(gnd),
	.combout(\ramstore~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~2 .lut_mask = 16'hF3C0;
defparam \ramstore~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N22
cycloneive_lcell_comb \ramstore~3 (
// Equation(s):
// \ramstore~3_combout  = (\syif.tbCTRL~input_o  & (\syif.store[3]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_3)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[3]~input_o ),
	.datad(\CPU|DP|rdata2_M [3]),
	.cin(gnd),
	.combout(\ramstore~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~3 .lut_mask = 16'hF3C0;
defparam \ramstore~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N22
cycloneive_lcell_comb \ramstore~4 (
// Equation(s):
// \ramstore~4_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[4]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_4))

	.dataa(\CPU|DP|rdata2_M [4]),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.store[4]~input_o ),
	.cin(gnd),
	.combout(\ramstore~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~4 .lut_mask = 16'hFA0A;
defparam \ramstore~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N24
cycloneive_lcell_comb \ramstore~5 (
// Equation(s):
// \ramstore~5_combout  = (\syif.tbCTRL~input_o  & (\syif.store[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_5)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[5]~input_o ),
	.datad(\CPU|DP|rdata2_M [5]),
	.cin(gnd),
	.combout(\ramstore~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~5 .lut_mask = 16'hF3C0;
defparam \ramstore~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N22
cycloneive_lcell_comb \ramstore~6 (
// Equation(s):
// \ramstore~6_combout  = (\syif.tbCTRL~input_o  & (\syif.store[6]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_6)))

	.dataa(\syif.store[6]~input_o ),
	.datab(\CPU|DP|rdata2_M [6]),
	.datac(gnd),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~6 .lut_mask = 16'hAACC;
defparam \ramstore~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N0
cycloneive_lcell_comb \ramstore~7 (
// Equation(s):
// \ramstore~7_combout  = (\syif.tbCTRL~input_o  & (\syif.store[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_7)))

	.dataa(gnd),
	.datab(\syif.store[7]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rdata2_M [7]),
	.cin(gnd),
	.combout(\ramstore~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~7 .lut_mask = 16'hCFC0;
defparam \ramstore~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N22
cycloneive_lcell_comb \ramstore~8 (
// Equation(s):
// \ramstore~8_combout  = (\syif.tbCTRL~input_o  & (\syif.store[8]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_8)))

	.dataa(\syif.store[8]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rdata2_M [8]),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramstore~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~8 .lut_mask = 16'hB8B8;
defparam \ramstore~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N8
cycloneive_lcell_comb \ramstore~9 (
// Equation(s):
// \ramstore~9_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[9]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_9))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rdata2_M [9]),
	.datad(\syif.store[9]~input_o ),
	.cin(gnd),
	.combout(\ramstore~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~9 .lut_mask = 16'hFC30;
defparam \ramstore~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N22
cycloneive_lcell_comb \ramstore~10 (
// Equation(s):
// \ramstore~10_combout  = (\syif.tbCTRL~input_o  & (\syif.store[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_10)))

	.dataa(\syif.store[10]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rdata2_M [10]),
	.cin(gnd),
	.combout(\ramstore~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~10 .lut_mask = 16'hAFA0;
defparam \ramstore~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N26
cycloneive_lcell_comb \ramstore~11 (
// Equation(s):
// \ramstore~11_combout  = (\syif.tbCTRL~input_o  & (\syif.store[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_11)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[11]~input_o ),
	.datad(\CPU|DP|rdata2_M [11]),
	.cin(gnd),
	.combout(\ramstore~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~11 .lut_mask = 16'hF3C0;
defparam \ramstore~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N18
cycloneive_lcell_comb \ramstore~12 (
// Equation(s):
// \ramstore~12_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[12]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_12))

	.dataa(\CPU|DP|rdata2_M [12]),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.store[12]~input_o ),
	.cin(gnd),
	.combout(\ramstore~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~12 .lut_mask = 16'hFA0A;
defparam \ramstore~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N16
cycloneive_lcell_comb \ramstore~13 (
// Equation(s):
// \ramstore~13_combout  = (\syif.tbCTRL~input_o  & (\syif.store[13]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_13)))

	.dataa(\syif.store[13]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rdata2_M [13]),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramstore~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~13 .lut_mask = 16'hB8B8;
defparam \ramstore~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N18
cycloneive_lcell_comb \ramstore~14 (
// Equation(s):
// \ramstore~14_combout  = (\syif.tbCTRL~input_o  & (\syif.store[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_14)))

	.dataa(\syif.store[14]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rdata2_M [14]),
	.cin(gnd),
	.combout(\ramstore~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~14 .lut_mask = 16'hAFA0;
defparam \ramstore~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N8
cycloneive_lcell_comb \ramstore~15 (
// Equation(s):
// \ramstore~15_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[15]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_15))

	.dataa(gnd),
	.datab(\CPU|DP|rdata2_M [15]),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.store[15]~input_o ),
	.cin(gnd),
	.combout(\ramstore~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~15 .lut_mask = 16'hFC0C;
defparam \ramstore~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N20
cycloneive_lcell_comb \ramstore~16 (
// Equation(s):
// \ramstore~16_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[16]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_16))

	.dataa(\CPU|DP|rdata2_M [16]),
	.datab(gnd),
	.datac(\syif.store[16]~input_o ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~16 .lut_mask = 16'hF0AA;
defparam \ramstore~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N4
cycloneive_lcell_comb \ramstore~17 (
// Equation(s):
// \ramstore~17_combout  = (\syif.tbCTRL~input_o  & (\syif.store[17]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_17)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[17]~input_o ),
	.datad(\CPU|DP|rdata2_M [17]),
	.cin(gnd),
	.combout(\ramstore~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~17 .lut_mask = 16'hF3C0;
defparam \ramstore~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N2
cycloneive_lcell_comb \ramstore~18 (
// Equation(s):
// \ramstore~18_combout  = (\syif.tbCTRL~input_o  & (\syif.store[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_18)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[18]~input_o ),
	.datad(\CPU|DP|rdata2_M [18]),
	.cin(gnd),
	.combout(\ramstore~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~18 .lut_mask = 16'hF3C0;
defparam \ramstore~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N18
cycloneive_lcell_comb \ramstore~19 (
// Equation(s):
// \ramstore~19_combout  = (\syif.tbCTRL~input_o  & (\syif.store[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_19)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[19]~input_o ),
	.datad(\CPU|DP|rdata2_M [19]),
	.cin(gnd),
	.combout(\ramstore~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~19 .lut_mask = 16'hF3C0;
defparam \ramstore~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N20
cycloneive_lcell_comb \ramstore~20 (
// Equation(s):
// \ramstore~20_combout  = (\syif.tbCTRL~input_o  & (\syif.store[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_20)))

	.dataa(\syif.store[20]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rdata2_M [20]),
	.cin(gnd),
	.combout(\ramstore~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~20 .lut_mask = 16'hAFA0;
defparam \ramstore~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N8
cycloneive_lcell_comb \ramstore~21 (
// Equation(s):
// \ramstore~21_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[21]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_21))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|rdata2_M [21]),
	.datac(gnd),
	.datad(\syif.store[21]~input_o ),
	.cin(gnd),
	.combout(\ramstore~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~21 .lut_mask = 16'hEE44;
defparam \ramstore~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N30
cycloneive_lcell_comb \ramstore~22 (
// Equation(s):
// \ramstore~22_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[22]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_22))

	.dataa(\CPU|DP|rdata2_M [22]),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.store[22]~input_o ),
	.cin(gnd),
	.combout(\ramstore~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~22 .lut_mask = 16'hFA0A;
defparam \ramstore~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N16
cycloneive_lcell_comb \ramstore~23 (
// Equation(s):
// \ramstore~23_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[23]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_23))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|rdata2_M [23]),
	.datac(gnd),
	.datad(\syif.store[23]~input_o ),
	.cin(gnd),
	.combout(\ramstore~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~23 .lut_mask = 16'hEE44;
defparam \ramstore~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N30
cycloneive_lcell_comb \ramstore~24 (
// Equation(s):
// \ramstore~24_combout  = (\syif.tbCTRL~input_o  & (\syif.store[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_24)))

	.dataa(\syif.store[24]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rdata2_M [24]),
	.cin(gnd),
	.combout(\ramstore~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~24 .lut_mask = 16'hAFA0;
defparam \ramstore~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N28
cycloneive_lcell_comb \ramstore~25 (
// Equation(s):
// \ramstore~25_combout  = (\syif.tbCTRL~input_o  & (\syif.store[25]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_25)))

	.dataa(\syif.store[25]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|rdata2_M [25]),
	.cin(gnd),
	.combout(\ramstore~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~25 .lut_mask = 16'hBB88;
defparam \ramstore~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N8
cycloneive_lcell_comb \ramstore~26 (
// Equation(s):
// \ramstore~26_combout  = (\syif.tbCTRL~input_o  & (\syif.store[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_26)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[26]~input_o ),
	.datad(\CPU|DP|rdata2_M [26]),
	.cin(gnd),
	.combout(\ramstore~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~26 .lut_mask = 16'hF3C0;
defparam \ramstore~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N26
cycloneive_lcell_comb \ramstore~27 (
// Equation(s):
// \ramstore~27_combout  = (\syif.tbCTRL~input_o  & (\syif.store[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_27)))

	.dataa(gnd),
	.datab(\syif.store[27]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rdata2_M [27]),
	.cin(gnd),
	.combout(\ramstore~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~27 .lut_mask = 16'hCFC0;
defparam \ramstore~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N24
cycloneive_lcell_comb \ramstore~28 (
// Equation(s):
// \ramstore~28_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[28]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_28))

	.dataa(\CPU|DP|rdata2_M [28]),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.store[28]~input_o ),
	.cin(gnd),
	.combout(\ramstore~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~28 .lut_mask = 16'hFA0A;
defparam \ramstore~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N16
cycloneive_lcell_comb \ramstore~29 (
// Equation(s):
// \ramstore~29_combout  = (\syif.tbCTRL~input_o  & (\syif.store[29]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_29)))

	.dataa(\syif.store[29]~input_o ),
	.datab(gnd),
	.datac(\CPU|DP|rdata2_M [29]),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~29 .lut_mask = 16'hAAF0;
defparam \ramstore~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N4
cycloneive_lcell_comb \ramstore~30 (
// Equation(s):
// \ramstore~30_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[30]~input_o ))) # (!\syif.tbCTRL~input_o  & (rdata2_M_30))

	.dataa(gnd),
	.datab(\CPU|DP|rdata2_M [30]),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.store[30]~input_o ),
	.cin(gnd),
	.combout(\ramstore~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~30 .lut_mask = 16'hFC0C;
defparam \ramstore~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N14
cycloneive_lcell_comb \ramstore~31 (
// Equation(s):
// \ramstore~31_combout  = (\syif.tbCTRL~input_o  & (\syif.store[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((rdata2_M_31)))

	.dataa(gnd),
	.datab(\syif.store[31]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rdata2_M [31]),
	.cin(gnd),
	.combout(\ramstore~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~31 .lut_mask = 16'hCFC0;
defparam \ramstore~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N22
cycloneive_lcell_comb \ramaddr~29_wirecell (
// Equation(s):
// \ramaddr~29_wirecell_combout  = !\ramaddr~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\ramaddr~29_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29_wirecell .lut_mask = 16'h00FF;
defparam \ramaddr~29_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: JTAG_X1_Y37_N0
cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

// Location: FF_X45_Y33_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y32_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hA50A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .lut_mask = 16'hA5A5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X46_Y34_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y34_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y34_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y34_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y34_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y32_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .lut_mask = 16'hFC22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(gnd),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .lut_mask = 16'hF5A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .lut_mask = 16'hF4A4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .lut_mask = 16'hF1A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .lut_mask = 16'hAA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .lut_mask = 16'hBF80;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .lut_mask = 16'h002A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .lut_mask = 16'hBA88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .lut_mask = 16'hDC10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .lut_mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .lut_mask = 16'hC001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .lut_mask = 16'h0100;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .lut_mask = 16'hFF08;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .lut_mask = 16'h00F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .lut_mask = 16'h2A24;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .lut_mask = 16'hD2F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y33_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .lut_mask = 16'hBA10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .lut_mask = 16'hF0F1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .lut_mask = 16'h0100;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y33_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .lut_mask = 16'hFF20;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .lut_mask = 16'h5050;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .lut_mask = 16'h0054;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .lut_mask = 16'h0E0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .lut_mask = 16'hEEEC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .lut_mask = 16'hD5C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hFF20;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .lut_mask = 16'h3F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .lut_mask = 16'h23A8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 .lut_mask = 16'h001A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .lut_mask = 16'hE2E2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .lut_mask = 16'h138D;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .lut_mask = 16'h2A0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N8
cycloneive_io_ibuf \syif.addr[1]~input (
	.i(\syif.addr [1]),
	.ibar(gnd),
	.o(\syif.addr[1]~input_o ));
// synopsys translate_off
defparam \syif.addr[1]~input .bus_hold = "false";
defparam \syif.addr[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N1
cycloneive_io_ibuf \syif.tbCTRL~input (
	.i(\syif.tbCTRL ),
	.ibar(gnd),
	.o(\syif.tbCTRL~input_o ));
// synopsys translate_off
defparam \syif.tbCTRL~input .bus_hold = "false";
defparam \syif.tbCTRL~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y35_N22
cycloneive_io_ibuf \syif.addr[0]~input (
	.i(\syif.addr [0]),
	.ibar(gnd),
	.o(\syif.addr[0]~input_o ));
// synopsys translate_off
defparam \syif.addr[0]~input .bus_hold = "false";
defparam \syif.addr[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X38_Y73_N22
cycloneive_io_ibuf \syif.addr[3]~input (
	.i(\syif.addr [3]),
	.ibar(gnd),
	.o(\syif.addr[3]~input_o ));
// synopsys translate_off
defparam \syif.addr[3]~input .bus_hold = "false";
defparam \syif.addr[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y40_N8
cycloneive_io_ibuf \syif.addr[2]~input (
	.i(\syif.addr [2]),
	.ibar(gnd),
	.o(\syif.addr[2]~input_o ));
// synopsys translate_off
defparam \syif.addr[2]~input .bus_hold = "false";
defparam \syif.addr[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N1
cycloneive_io_ibuf \syif.addr[5]~input (
	.i(\syif.addr [5]),
	.ibar(gnd),
	.o(\syif.addr[5]~input_o ));
// synopsys translate_off
defparam \syif.addr[5]~input .bus_hold = "false";
defparam \syif.addr[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N15
cycloneive_io_ibuf \syif.addr[4]~input (
	.i(\syif.addr [4]),
	.ibar(gnd),
	.o(\syif.addr[4]~input_o ));
// synopsys translate_off
defparam \syif.addr[4]~input .bus_hold = "false";
defparam \syif.addr[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N1
cycloneive_io_ibuf \syif.addr[7]~input (
	.i(\syif.addr [7]),
	.ibar(gnd),
	.o(\syif.addr[7]~input_o ));
// synopsys translate_off
defparam \syif.addr[7]~input .bus_hold = "false";
defparam \syif.addr[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N8
cycloneive_io_ibuf \syif.addr[6]~input (
	.i(\syif.addr [6]),
	.ibar(gnd),
	.o(\syif.addr[6]~input_o ));
// synopsys translate_off
defparam \syif.addr[6]~input .bus_hold = "false";
defparam \syif.addr[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N8
cycloneive_io_ibuf \syif.addr[9]~input (
	.i(\syif.addr [9]),
	.ibar(gnd),
	.o(\syif.addr[9]~input_o ));
// synopsys translate_off
defparam \syif.addr[9]~input .bus_hold = "false";
defparam \syif.addr[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N15
cycloneive_io_ibuf \syif.addr[8]~input (
	.i(\syif.addr [8]),
	.ibar(gnd),
	.o(\syif.addr[8]~input_o ));
// synopsys translate_off
defparam \syif.addr[8]~input .bus_hold = "false";
defparam \syif.addr[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y73_N1
cycloneive_io_ibuf \syif.addr[11]~input (
	.i(\syif.addr [11]),
	.ibar(gnd),
	.o(\syif.addr[11]~input_o ));
// synopsys translate_off
defparam \syif.addr[11]~input .bus_hold = "false";
defparam \syif.addr[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N22
cycloneive_io_ibuf \syif.addr[10]~input (
	.i(\syif.addr [10]),
	.ibar(gnd),
	.o(\syif.addr[10]~input_o ));
// synopsys translate_off
defparam \syif.addr[10]~input .bus_hold = "false";
defparam \syif.addr[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N22
cycloneive_io_ibuf \syif.addr[13]~input (
	.i(\syif.addr [13]),
	.ibar(gnd),
	.o(\syif.addr[13]~input_o ));
// synopsys translate_off
defparam \syif.addr[13]~input .bus_hold = "false";
defparam \syif.addr[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y40_N1
cycloneive_io_ibuf \syif.addr[12]~input (
	.i(\syif.addr [12]),
	.ibar(gnd),
	.o(\syif.addr[12]~input_o ));
// synopsys translate_off
defparam \syif.addr[12]~input .bus_hold = "false";
defparam \syif.addr[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N15
cycloneive_io_ibuf \syif.addr[15]~input (
	.i(\syif.addr [15]),
	.ibar(gnd),
	.o(\syif.addr[15]~input_o ));
// synopsys translate_off
defparam \syif.addr[15]~input .bus_hold = "false";
defparam \syif.addr[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y73_N8
cycloneive_io_ibuf \syif.addr[14]~input (
	.i(\syif.addr [14]),
	.ibar(gnd),
	.o(\syif.addr[14]~input_o ));
// synopsys translate_off
defparam \syif.addr[14]~input .bus_hold = "false";
defparam \syif.addr[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N1
cycloneive_io_ibuf \syif.addr[17]~input (
	.i(\syif.addr [17]),
	.ibar(gnd),
	.o(\syif.addr[17]~input_o ));
// synopsys translate_off
defparam \syif.addr[17]~input .bus_hold = "false";
defparam \syif.addr[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y73_N8
cycloneive_io_ibuf \syif.addr[16]~input (
	.i(\syif.addr [16]),
	.ibar(gnd),
	.o(\syif.addr[16]~input_o ));
// synopsys translate_off
defparam \syif.addr[16]~input .bus_hold = "false";
defparam \syif.addr[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N15
cycloneive_io_ibuf \syif.addr[19]~input (
	.i(\syif.addr [19]),
	.ibar(gnd),
	.o(\syif.addr[19]~input_o ));
// synopsys translate_off
defparam \syif.addr[19]~input .bus_hold = "false";
defparam \syif.addr[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N8
cycloneive_io_ibuf \syif.addr[18]~input (
	.i(\syif.addr [18]),
	.ibar(gnd),
	.o(\syif.addr[18]~input_o ));
// synopsys translate_off
defparam \syif.addr[18]~input .bus_hold = "false";
defparam \syif.addr[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N22
cycloneive_io_ibuf \syif.addr[21]~input (
	.i(\syif.addr [21]),
	.ibar(gnd),
	.o(\syif.addr[21]~input_o ));
// synopsys translate_off
defparam \syif.addr[21]~input .bus_hold = "false";
defparam \syif.addr[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N22
cycloneive_io_ibuf \syif.addr[20]~input (
	.i(\syif.addr [20]),
	.ibar(gnd),
	.o(\syif.addr[20]~input_o ));
// synopsys translate_off
defparam \syif.addr[20]~input .bus_hold = "false";
defparam \syif.addr[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N15
cycloneive_io_ibuf \syif.addr[23]~input (
	.i(\syif.addr [23]),
	.ibar(gnd),
	.o(\syif.addr[23]~input_o ));
// synopsys translate_off
defparam \syif.addr[23]~input .bus_hold = "false";
defparam \syif.addr[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N8
cycloneive_io_ibuf \syif.addr[22]~input (
	.i(\syif.addr [22]),
	.ibar(gnd),
	.o(\syif.addr[22]~input_o ));
// synopsys translate_off
defparam \syif.addr[22]~input .bus_hold = "false";
defparam \syif.addr[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N1
cycloneive_io_ibuf \syif.addr[25]~input (
	.i(\syif.addr [25]),
	.ibar(gnd),
	.o(\syif.addr[25]~input_o ));
// synopsys translate_off
defparam \syif.addr[25]~input .bus_hold = "false";
defparam \syif.addr[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N1
cycloneive_io_ibuf \syif.addr[24]~input (
	.i(\syif.addr [24]),
	.ibar(gnd),
	.o(\syif.addr[24]~input_o ));
// synopsys translate_off
defparam \syif.addr[24]~input .bus_hold = "false";
defparam \syif.addr[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N15
cycloneive_io_ibuf \syif.addr[27]~input (
	.i(\syif.addr [27]),
	.ibar(gnd),
	.o(\syif.addr[27]~input_o ));
// synopsys translate_off
defparam \syif.addr[27]~input .bus_hold = "false";
defparam \syif.addr[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N15
cycloneive_io_ibuf \syif.addr[26]~input (
	.i(\syif.addr [26]),
	.ibar(gnd),
	.o(\syif.addr[26]~input_o ));
// synopsys translate_off
defparam \syif.addr[26]~input .bus_hold = "false";
defparam \syif.addr[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N1
cycloneive_io_ibuf \syif.addr[29]~input (
	.i(\syif.addr [29]),
	.ibar(gnd),
	.o(\syif.addr[29]~input_o ));
// synopsys translate_off
defparam \syif.addr[29]~input .bus_hold = "false";
defparam \syif.addr[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N8
cycloneive_io_ibuf \syif.addr[28]~input (
	.i(\syif.addr [28]),
	.ibar(gnd),
	.o(\syif.addr[28]~input_o ));
// synopsys translate_off
defparam \syif.addr[28]~input .bus_hold = "false";
defparam \syif.addr[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y73_N8
cycloneive_io_ibuf \syif.addr[31]~input (
	.i(\syif.addr [31]),
	.ibar(gnd),
	.o(\syif.addr[31]~input_o ));
// synopsys translate_off
defparam \syif.addr[31]~input .bus_hold = "false";
defparam \syif.addr[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N15
cycloneive_io_ibuf \syif.addr[30]~input (
	.i(\syif.addr [30]),
	.ibar(gnd),
	.o(\syif.addr[30]~input_o ));
// synopsys translate_off
defparam \syif.addr[30]~input .bus_hold = "false";
defparam \syif.addr[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y73_N1
cycloneive_io_ibuf \syif.WEN~input (
	.i(\syif.WEN ),
	.ibar(gnd),
	.o(\syif.WEN~input_o ));
// synopsys translate_off
defparam \syif.WEN~input .bus_hold = "false";
defparam \syif.WEN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N22
cycloneive_io_ibuf \syif.REN~input (
	.i(\syif.REN ),
	.ibar(gnd),
	.o(\syif.REN~input_o ));
// synopsys translate_off
defparam \syif.REN~input .bus_hold = "false";
defparam \syif.REN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N15
cycloneive_io_ibuf \nRST~input (
	.i(nRST),
	.ibar(gnd),
	.o(\nRST~input_o ));
// synopsys translate_off
defparam \nRST~input .bus_hold = "false";
defparam \nRST~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N8
cycloneive_io_ibuf \CLK~input (
	.i(CLK),
	.ibar(gnd),
	.o(\CLK~input_o ));
// synopsys translate_off
defparam \CLK~input .bus_hold = "false";
defparam \CLK~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y33_N8
cycloneive_io_ibuf \syif.store[0]~input (
	.i(\syif.store [0]),
	.ibar(gnd),
	.o(\syif.store[0]~input_o ));
// synopsys translate_off
defparam \syif.store[0]~input .bus_hold = "false";
defparam \syif.store[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N22
cycloneive_io_ibuf \syif.store[1]~input (
	.i(\syif.store [1]),
	.ibar(gnd),
	.o(\syif.store[1]~input_o ));
// synopsys translate_off
defparam \syif.store[1]~input .bus_hold = "false";
defparam \syif.store[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N22
cycloneive_io_ibuf \syif.store[2]~input (
	.i(\syif.store [2]),
	.ibar(gnd),
	.o(\syif.store[2]~input_o ));
// synopsys translate_off
defparam \syif.store[2]~input .bus_hold = "false";
defparam \syif.store[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y73_N22
cycloneive_io_ibuf \syif.store[3]~input (
	.i(\syif.store [3]),
	.ibar(gnd),
	.o(\syif.store[3]~input_o ));
// synopsys translate_off
defparam \syif.store[3]~input .bus_hold = "false";
defparam \syif.store[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y73_N8
cycloneive_io_ibuf \syif.store[4]~input (
	.i(\syif.store [4]),
	.ibar(gnd),
	.o(\syif.store[4]~input_o ));
// synopsys translate_off
defparam \syif.store[4]~input .bus_hold = "false";
defparam \syif.store[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y73_N15
cycloneive_io_ibuf \syif.store[5]~input (
	.i(\syif.store [5]),
	.ibar(gnd),
	.o(\syif.store[5]~input_o ));
// synopsys translate_off
defparam \syif.store[5]~input .bus_hold = "false";
defparam \syif.store[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y73_N22
cycloneive_io_ibuf \syif.store[6]~input (
	.i(\syif.store [6]),
	.ibar(gnd),
	.o(\syif.store[6]~input_o ));
// synopsys translate_off
defparam \syif.store[6]~input .bus_hold = "false";
defparam \syif.store[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N1
cycloneive_io_ibuf \syif.store[7]~input (
	.i(\syif.store [7]),
	.ibar(gnd),
	.o(\syif.store[7]~input_o ));
// synopsys translate_off
defparam \syif.store[7]~input .bus_hold = "false";
defparam \syif.store[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N8
cycloneive_io_ibuf \syif.store[8]~input (
	.i(\syif.store [8]),
	.ibar(gnd),
	.o(\syif.store[8]~input_o ));
// synopsys translate_off
defparam \syif.store[8]~input .bus_hold = "false";
defparam \syif.store[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N8
cycloneive_io_ibuf \syif.store[9]~input (
	.i(\syif.store [9]),
	.ibar(gnd),
	.o(\syif.store[9]~input_o ));
// synopsys translate_off
defparam \syif.store[9]~input .bus_hold = "false";
defparam \syif.store[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N1
cycloneive_io_ibuf \syif.store[10]~input (
	.i(\syif.store [10]),
	.ibar(gnd),
	.o(\syif.store[10]~input_o ));
// synopsys translate_off
defparam \syif.store[10]~input .bus_hold = "false";
defparam \syif.store[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N1
cycloneive_io_ibuf \syif.store[11]~input (
	.i(\syif.store [11]),
	.ibar(gnd),
	.o(\syif.store[11]~input_o ));
// synopsys translate_off
defparam \syif.store[11]~input .bus_hold = "false";
defparam \syif.store[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N1
cycloneive_io_ibuf \syif.store[12]~input (
	.i(\syif.store [12]),
	.ibar(gnd),
	.o(\syif.store[12]~input_o ));
// synopsys translate_off
defparam \syif.store[12]~input .bus_hold = "false";
defparam \syif.store[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y73_N1
cycloneive_io_ibuf \syif.store[13]~input (
	.i(\syif.store [13]),
	.ibar(gnd),
	.o(\syif.store[13]~input_o ));
// synopsys translate_off
defparam \syif.store[13]~input .bus_hold = "false";
defparam \syif.store[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y33_N1
cycloneive_io_ibuf \syif.store[14]~input (
	.i(\syif.store [14]),
	.ibar(gnd),
	.o(\syif.store[14]~input_o ));
// synopsys translate_off
defparam \syif.store[14]~input .bus_hold = "false";
defparam \syif.store[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N22
cycloneive_io_ibuf \syif.store[15]~input (
	.i(\syif.store [15]),
	.ibar(gnd),
	.o(\syif.store[15]~input_o ));
// synopsys translate_off
defparam \syif.store[15]~input .bus_hold = "false";
defparam \syif.store[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N15
cycloneive_io_ibuf \syif.store[16]~input (
	.i(\syif.store [16]),
	.ibar(gnd),
	.o(\syif.store[16]~input_o ));
// synopsys translate_off
defparam \syif.store[16]~input .bus_hold = "false";
defparam \syif.store[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y32_N8
cycloneive_io_ibuf \syif.store[17]~input (
	.i(\syif.store [17]),
	.ibar(gnd),
	.o(\syif.store[17]~input_o ));
// synopsys translate_off
defparam \syif.store[17]~input .bus_hold = "false";
defparam \syif.store[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y31_N8
cycloneive_io_ibuf \syif.store[18]~input (
	.i(\syif.store [18]),
	.ibar(gnd),
	.o(\syif.store[18]~input_o ));
// synopsys translate_off
defparam \syif.store[18]~input .bus_hold = "false";
defparam \syif.store[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N8
cycloneive_io_ibuf \syif.store[19]~input (
	.i(\syif.store [19]),
	.ibar(gnd),
	.o(\syif.store[19]~input_o ));
// synopsys translate_off
defparam \syif.store[19]~input .bus_hold = "false";
defparam \syif.store[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X81_Y73_N22
cycloneive_io_ibuf \syif.store[20]~input (
	.i(\syif.store [20]),
	.ibar(gnd),
	.o(\syif.store[20]~input_o ));
// synopsys translate_off
defparam \syif.store[20]~input .bus_hold = "false";
defparam \syif.store[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N1
cycloneive_io_ibuf \syif.store[21]~input (
	.i(\syif.store [21]),
	.ibar(gnd),
	.o(\syif.store[21]~input_o ));
// synopsys translate_off
defparam \syif.store[21]~input .bus_hold = "false";
defparam \syif.store[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y73_N22
cycloneive_io_ibuf \syif.store[22]~input (
	.i(\syif.store [22]),
	.ibar(gnd),
	.o(\syif.store[22]~input_o ));
// synopsys translate_off
defparam \syif.store[22]~input .bus_hold = "false";
defparam \syif.store[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N15
cycloneive_io_ibuf \syif.store[23]~input (
	.i(\syif.store [23]),
	.ibar(gnd),
	.o(\syif.store[23]~input_o ));
// synopsys translate_off
defparam \syif.store[23]~input .bus_hold = "false";
defparam \syif.store[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y73_N15
cycloneive_io_ibuf \syif.store[24]~input (
	.i(\syif.store [24]),
	.ibar(gnd),
	.o(\syif.store[24]~input_o ));
// synopsys translate_off
defparam \syif.store[24]~input .bus_hold = "false";
defparam \syif.store[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N8
cycloneive_io_ibuf \syif.store[25]~input (
	.i(\syif.store [25]),
	.ibar(gnd),
	.o(\syif.store[25]~input_o ));
// synopsys translate_off
defparam \syif.store[25]~input .bus_hold = "false";
defparam \syif.store[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N15
cycloneive_io_ibuf \syif.store[26]~input (
	.i(\syif.store [26]),
	.ibar(gnd),
	.o(\syif.store[26]~input_o ));
// synopsys translate_off
defparam \syif.store[26]~input .bus_hold = "false";
defparam \syif.store[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y73_N1
cycloneive_io_ibuf \syif.store[27]~input (
	.i(\syif.store [27]),
	.ibar(gnd),
	.o(\syif.store[27]~input_o ));
// synopsys translate_off
defparam \syif.store[27]~input .bus_hold = "false";
defparam \syif.store[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N1
cycloneive_io_ibuf \syif.store[28]~input (
	.i(\syif.store [28]),
	.ibar(gnd),
	.o(\syif.store[28]~input_o ));
// synopsys translate_off
defparam \syif.store[28]~input .bus_hold = "false";
defparam \syif.store[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N8
cycloneive_io_ibuf \syif.store[29]~input (
	.i(\syif.store [29]),
	.ibar(gnd),
	.o(\syif.store[29]~input_o ));
// synopsys translate_off
defparam \syif.store[29]~input .bus_hold = "false";
defparam \syif.store[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y41_N1
cycloneive_io_ibuf \syif.store[30]~input (
	.i(\syif.store [30]),
	.ibar(gnd),
	.o(\syif.store[30]~input_o ));
// synopsys translate_off
defparam \syif.store[30]~input .bus_hold = "false";
defparam \syif.store[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N1
cycloneive_io_ibuf \syif.store[31]~input (
	.i(\syif.store [31]),
	.ibar(gnd),
	.o(\syif.store[31]~input_o ));
// synopsys translate_off
defparam \syif.store[31]~input .bus_hold = "false";
defparam \syif.store[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G4
cycloneive_clkctrl \nRST~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\nRST~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\nRST~inputclkctrl_outclk ));
// synopsys translate_off
defparam \nRST~inputclkctrl .clock_type = "global clock";
defparam \nRST~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G3
cycloneive_clkctrl \altera_internal_jtag~TCKUTAPclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\altera_internal_jtag~TCKUTAP }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ));
// synopsys translate_off
defparam \altera_internal_jtag~TCKUTAPclkctrl .clock_type = "global clock";
defparam \altera_internal_jtag~TCKUTAPclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G2
cycloneive_clkctrl \CLK~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CLK~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CLK~inputclkctrl_outclk ));
// synopsys translate_off
defparam \CLK~inputclkctrl .clock_type = "global clock";
defparam \CLK~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N9
cycloneive_io_obuf \syif.halt~output (
	.i(\CPU|DP|halt_WB~q ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.halt ),
	.obar());
// synopsys translate_off
defparam \syif.halt~output .bus_hold = "false";
defparam \syif.halt~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y31_N2
cycloneive_io_obuf \syif.load[0]~output (
	.i(\RAM|ramif.ramload[0]~0_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [0]),
	.obar());
// synopsys translate_off
defparam \syif.load[0]~output .bus_hold = "false";
defparam \syif.load[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N2
cycloneive_io_obuf \syif.load[1]~output (
	.i(\RAM|ramif.ramload[1]~1_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [1]),
	.obar());
// synopsys translate_off
defparam \syif.load[1]~output .bus_hold = "false";
defparam \syif.load[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y0_N23
cycloneive_io_obuf \syif.load[2]~output (
	.i(\RAM|ramif.ramload[2]~2_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [2]),
	.obar());
// synopsys translate_off
defparam \syif.load[2]~output .bus_hold = "false";
defparam \syif.load[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N23
cycloneive_io_obuf \syif.load[3]~output (
	.i(\RAM|ramif.ramload[3]~3_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [3]),
	.obar());
// synopsys translate_off
defparam \syif.load[3]~output .bus_hold = "false";
defparam \syif.load[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y34_N16
cycloneive_io_obuf \syif.load[4]~output (
	.i(\RAM|ramif.ramload[4]~4_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [4]),
	.obar());
// synopsys translate_off
defparam \syif.load[4]~output .bus_hold = "false";
defparam \syif.load[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N2
cycloneive_io_obuf \syif.load[5]~output (
	.i(\RAM|ramif.ramload[5]~5_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [5]),
	.obar());
// synopsys translate_off
defparam \syif.load[5]~output .bus_hold = "false";
defparam \syif.load[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N16
cycloneive_io_obuf \syif.load[6]~output (
	.i(\RAM|ramif.ramload[6]~6_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [6]),
	.obar());
// synopsys translate_off
defparam \syif.load[6]~output .bus_hold = "false";
defparam \syif.load[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y73_N16
cycloneive_io_obuf \syif.load[7]~output (
	.i(\RAM|ramif.ramload[7]~7_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [7]),
	.obar());
// synopsys translate_off
defparam \syif.load[7]~output .bus_hold = "false";
defparam \syif.load[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y73_N23
cycloneive_io_obuf \syif.load[8]~output (
	.i(\RAM|ramif.ramload[8]~8_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [8]),
	.obar());
// synopsys translate_off
defparam \syif.load[8]~output .bus_hold = "false";
defparam \syif.load[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N2
cycloneive_io_obuf \syif.load[9]~output (
	.i(\RAM|ramif.ramload[9]~9_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [9]),
	.obar());
// synopsys translate_off
defparam \syif.load[9]~output .bus_hold = "false";
defparam \syif.load[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N23
cycloneive_io_obuf \syif.load[10]~output (
	.i(\RAM|ramif.ramload[10]~10_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [10]),
	.obar());
// synopsys translate_off
defparam \syif.load[10]~output .bus_hold = "false";
defparam \syif.load[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N9
cycloneive_io_obuf \syif.load[11]~output (
	.i(\RAM|ramif.ramload[11]~11_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [11]),
	.obar());
// synopsys translate_off
defparam \syif.load[11]~output .bus_hold = "false";
defparam \syif.load[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y73_N16
cycloneive_io_obuf \syif.load[12]~output (
	.i(\RAM|ramif.ramload[12]~12_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [12]),
	.obar());
// synopsys translate_off
defparam \syif.load[12]~output .bus_hold = "false";
defparam \syif.load[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X69_Y73_N16
cycloneive_io_obuf \syif.load[13]~output (
	.i(\RAM|ramif.ramload[13]~13_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [13]),
	.obar());
// synopsys translate_off
defparam \syif.load[13]~output .bus_hold = "false";
defparam \syif.load[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N16
cycloneive_io_obuf \syif.load[14]~output (
	.i(\RAM|ramif.ramload[14]~14_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [14]),
	.obar());
// synopsys translate_off
defparam \syif.load[14]~output .bus_hold = "false";
defparam \syif.load[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N2
cycloneive_io_obuf \syif.load[15]~output (
	.i(\RAM|ramif.ramload[15]~15_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [15]),
	.obar());
// synopsys translate_off
defparam \syif.load[15]~output .bus_hold = "false";
defparam \syif.load[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X79_Y73_N9
cycloneive_io_obuf \syif.load[16]~output (
	.i(\RAM|ramif.ramload[16]~16_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [16]),
	.obar());
// synopsys translate_off
defparam \syif.load[16]~output .bus_hold = "false";
defparam \syif.load[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y73_N9
cycloneive_io_obuf \syif.load[17]~output (
	.i(\RAM|ramif.ramload[17]~17_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [17]),
	.obar());
// synopsys translate_off
defparam \syif.load[17]~output .bus_hold = "false";
defparam \syif.load[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y35_N16
cycloneive_io_obuf \syif.load[18]~output (
	.i(\RAM|ramif.ramload[18]~18_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [18]),
	.obar());
// synopsys translate_off
defparam \syif.load[18]~output .bus_hold = "false";
defparam \syif.load[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X79_Y73_N2
cycloneive_io_obuf \syif.load[19]~output (
	.i(\RAM|ramif.ramload[19]~19_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [19]),
	.obar());
// synopsys translate_off
defparam \syif.load[19]~output .bus_hold = "false";
defparam \syif.load[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N9
cycloneive_io_obuf \syif.load[20]~output (
	.i(\RAM|ramif.ramload[20]~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [20]),
	.obar());
// synopsys translate_off
defparam \syif.load[20]~output .bus_hold = "false";
defparam \syif.load[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N23
cycloneive_io_obuf \syif.load[21]~output (
	.i(\RAM|ramif.ramload[21]~21_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [21]),
	.obar());
// synopsys translate_off
defparam \syif.load[21]~output .bus_hold = "false";
defparam \syif.load[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N23
cycloneive_io_obuf \syif.load[22]~output (
	.i(\RAM|ramif.ramload[22]~22_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [22]),
	.obar());
// synopsys translate_off
defparam \syif.load[22]~output .bus_hold = "false";
defparam \syif.load[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N2
cycloneive_io_obuf \syif.load[23]~output (
	.i(\RAM|ramif.ramload[23]~23_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [23]),
	.obar());
// synopsys translate_off
defparam \syif.load[23]~output .bus_hold = "false";
defparam \syif.load[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y73_N23
cycloneive_io_obuf \syif.load[24]~output (
	.i(\RAM|ramif.ramload[24]~24_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [24]),
	.obar());
// synopsys translate_off
defparam \syif.load[24]~output .bus_hold = "false";
defparam \syif.load[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N16
cycloneive_io_obuf \syif.load[25]~output (
	.i(\RAM|ramif.ramload[25]~25_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [25]),
	.obar());
// synopsys translate_off
defparam \syif.load[25]~output .bus_hold = "false";
defparam \syif.load[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N9
cycloneive_io_obuf \syif.load[26]~output (
	.i(\RAM|ramif.ramload[26]~26_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [26]),
	.obar());
// synopsys translate_off
defparam \syif.load[26]~output .bus_hold = "false";
defparam \syif.load[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N9
cycloneive_io_obuf \syif.load[27]~output (
	.i(\RAM|ramif.ramload[27]~27_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [27]),
	.obar());
// synopsys translate_off
defparam \syif.load[27]~output .bus_hold = "false";
defparam \syif.load[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N16
cycloneive_io_obuf \syif.load[28]~output (
	.i(\RAM|ramif.ramload[28]~28_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [28]),
	.obar());
// synopsys translate_off
defparam \syif.load[28]~output .bus_hold = "false";
defparam \syif.load[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N16
cycloneive_io_obuf \syif.load[29]~output (
	.i(\RAM|ramif.ramload[29]~29_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [29]),
	.obar());
// synopsys translate_off
defparam \syif.load[29]~output .bus_hold = "false";
defparam \syif.load[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y73_N9
cycloneive_io_obuf \syif.load[30]~output (
	.i(\RAM|ramif.ramload[30]~30_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [30]),
	.obar());
// synopsys translate_off
defparam \syif.load[30]~output .bus_hold = "false";
defparam \syif.load[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y32_N2
cycloneive_io_obuf \syif.load[31]~output (
	.i(\RAM|ramif.ramload[31]~31_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [31]),
	.obar());
// synopsys translate_off
defparam \syif.load[31]~output .bus_hold = "false";
defparam \syif.load[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y37_N1
cycloneive_io_obuf \altera_reserved_tdo~output (
	.i(\altera_internal_jtag~TDO ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(altera_reserved_tdo),
	.obar());
// synopsys translate_off
defparam \altera_reserved_tdo~output .bus_hold = "false";
defparam \altera_reserved_tdo~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOIBUF_X0_Y38_N1
cycloneive_io_ibuf \altera_reserved_tms~input (
	.i(altera_reserved_tms),
	.ibar(gnd),
	.o(\altera_reserved_tms~input_o ));
// synopsys translate_off
defparam \altera_reserved_tms~input .bus_hold = "false";
defparam \altera_reserved_tms~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y39_N1
cycloneive_io_ibuf \altera_reserved_tck~input (
	.i(altera_reserved_tck),
	.ibar(gnd),
	.o(\altera_reserved_tck~input_o ));
// synopsys translate_off
defparam \altera_reserved_tck~input .bus_hold = "false";
defparam \altera_reserved_tck~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y40_N1
cycloneive_io_ibuf \altera_reserved_tdi~input (
	.i(altera_reserved_tdi),
	.ibar(gnd),
	.o(\altera_reserved_tdi~input_o ));
// synopsys translate_off
defparam \altera_reserved_tdi~input .bus_hold = "false";
defparam \altera_reserved_tdi~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .lut_mask = 16'hFFFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .lut_mask = 16'hFFFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hE0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .lut_mask = 16'hF0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .lut_mask = 16'hFFFD;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .lut_mask = 16'hF0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y33_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .lut_mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N8
cycloneive_lcell_comb \~QIC_CREATED_GND~I (
// Equation(s):
// \~QIC_CREATED_GND~I_combout  = GND

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.cout());
// synopsys translate_off
defparam \~QIC_CREATED_GND~I .lut_mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .lut_mask = 16'hA080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .lut_mask = 16'h7430;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .lut_mask = 16'h0A0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .lut_mask = 16'h5AF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .lut_mask = 16'h5575;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .lut_mask = 16'h0001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .lut_mask = 16'h0010;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .lut_mask = 16'h1000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.asdata(\~QIC_CREATED_GND~I_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .lut_mask = 16'h00C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .lut_mask = 16'h7250;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .lut_mask = 16'hF0AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datac(gnd),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .lut_mask = 16'hCACA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .lut_mask = 16'hE040;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .lut_mask = 16'hCFC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y34_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .lut_mask = 16'hFA50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 (
	.dataa(gnd),
	.datab(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .lut_mask = 16'hCFC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 (
	.dataa(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .lut_mask = 16'hAFA0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .lut_mask = 16'h2000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .lut_mask = 16'h4400;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .lut_mask = 16'h1000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .lut_mask = 16'h55AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .lut_mask = 16'h0011;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .lut_mask = 16'hABAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16 .lut_mask = 16'hEAC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~10 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9 .lut_mask = 16'h3CCF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X43_Y32_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~10 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X43_Y32_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13 .lut_mask = 16'h3C3C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X43_Y32_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y32_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~11 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 .lut_mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .lut_mask = 16'hCCAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .lut_mask = 16'h010B;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .lut_mask = 16'h02E2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .lut_mask = 16'hCFC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .lut_mask = 16'hCCAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .lut_mask = 16'h6A54;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .lut_mask = 16'h3034;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .lut_mask = 16'hBB88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .lut_mask = 16'h3F3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .lut_mask = 16'hFAF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .lut_mask = 16'h07F5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo (
	.clk(!\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y36_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y59_N0
cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline (
	pc_out_3,
	pc_out_2,
	pc_out_5,
	pc_out_4,
	pc_out_7,
	pc_out_6,
	pc_out_9,
	pc_out_8,
	pc_out_11,
	pc_out_10,
	pc_out_13,
	pc_out_12,
	pc_out_15,
	pc_out_14,
	pc_out_17,
	pc_out_16,
	pc_out_19,
	pc_out_18,
	pc_out_21,
	pc_out_20,
	pc_out_23,
	pc_out_22,
	pc_out_25,
	pc_out_24,
	pc_out_27,
	pc_out_26,
	rdata2_M_0,
	rdata2_M_1,
	rdata2_M_2,
	rdata2_M_3,
	rdata2_M_4,
	rdata2_M_5,
	rdata2_M_6,
	rdata2_M_7,
	rdata2_M_8,
	rdata2_M_9,
	rdata2_M_10,
	rdata2_M_11,
	rdata2_M_12,
	rdata2_M_13,
	rdata2_M_14,
	rdata2_M_15,
	rdata2_M_16,
	rdata2_M_17,
	rdata2_M_18,
	rdata2_M_19,
	rdata2_M_20,
	rdata2_M_21,
	rdata2_M_22,
	rdata2_M_23,
	rdata2_M_24,
	rdata2_M_25,
	rdata2_M_26,
	rdata2_M_27,
	rdata2_M_28,
	rdata2_M_29,
	rdata2_M_30,
	rdata2_M_31,
	LessThan1,
	porto_M_1,
	pc_out_1,
	dWEN_M,
	dREN_M,
	porto_M_0,
	pc_out_0,
	porto_M_3,
	porto_M_2,
	porto_M_5,
	porto_M_4,
	porto_M_7,
	porto_M_6,
	porto_M_9,
	porto_M_8,
	porto_M_11,
	porto_M_10,
	porto_M_13,
	porto_M_12,
	porto_M_15,
	porto_M_14,
	porto_M_17,
	porto_M_16,
	porto_M_19,
	porto_M_18,
	porto_M_21,
	porto_M_20,
	porto_M_23,
	porto_M_22,
	porto_M_25,
	porto_M_24,
	porto_M_27,
	porto_M_26,
	porto_M_29,
	pc_out_29,
	porto_M_28,
	pc_out_28,
	porto_M_31,
	pc_out_31,
	porto_M_30,
	pc_out_30,
	always0,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	nRST,
	nRST1,
	CLK,
	halt_WB,
	devpor,
	devclrn,
	devoe);
output 	pc_out_3;
output 	pc_out_2;
output 	pc_out_5;
output 	pc_out_4;
output 	pc_out_7;
output 	pc_out_6;
output 	pc_out_9;
output 	pc_out_8;
output 	pc_out_11;
output 	pc_out_10;
output 	pc_out_13;
output 	pc_out_12;
output 	pc_out_15;
output 	pc_out_14;
output 	pc_out_17;
output 	pc_out_16;
output 	pc_out_19;
output 	pc_out_18;
output 	pc_out_21;
output 	pc_out_20;
output 	pc_out_23;
output 	pc_out_22;
output 	pc_out_25;
output 	pc_out_24;
output 	pc_out_27;
output 	pc_out_26;
output 	rdata2_M_0;
output 	rdata2_M_1;
output 	rdata2_M_2;
output 	rdata2_M_3;
output 	rdata2_M_4;
output 	rdata2_M_5;
output 	rdata2_M_6;
output 	rdata2_M_7;
output 	rdata2_M_8;
output 	rdata2_M_9;
output 	rdata2_M_10;
output 	rdata2_M_11;
output 	rdata2_M_12;
output 	rdata2_M_13;
output 	rdata2_M_14;
output 	rdata2_M_15;
output 	rdata2_M_16;
output 	rdata2_M_17;
output 	rdata2_M_18;
output 	rdata2_M_19;
output 	rdata2_M_20;
output 	rdata2_M_21;
output 	rdata2_M_22;
output 	rdata2_M_23;
output 	rdata2_M_24;
output 	rdata2_M_25;
output 	rdata2_M_26;
output 	rdata2_M_27;
output 	rdata2_M_28;
output 	rdata2_M_29;
output 	rdata2_M_30;
output 	rdata2_M_31;
input 	LessThan1;
output 	porto_M_1;
output 	pc_out_1;
output 	dWEN_M;
output 	dREN_M;
output 	porto_M_0;
output 	pc_out_0;
output 	porto_M_3;
output 	porto_M_2;
output 	porto_M_5;
output 	porto_M_4;
output 	porto_M_7;
output 	porto_M_6;
output 	porto_M_9;
output 	porto_M_8;
output 	porto_M_11;
output 	porto_M_10;
output 	porto_M_13;
output 	porto_M_12;
output 	porto_M_15;
output 	porto_M_14;
output 	porto_M_17;
output 	porto_M_16;
output 	porto_M_19;
output 	porto_M_18;
output 	porto_M_21;
output 	porto_M_20;
output 	porto_M_23;
output 	porto_M_22;
output 	porto_M_25;
output 	porto_M_24;
output 	porto_M_27;
output 	porto_M_26;
output 	porto_M_29;
output 	pc_out_29;
output 	porto_M_28;
output 	pc_out_28;
output 	porto_M_31;
output 	pc_out_31;
output 	porto_M_30;
output 	pc_out_30;
input 	always0;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	nRST;
input 	nRST1;
input 	CLK;
output 	halt_WB;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \CM|dhit~0_combout ;
wire \CC|iwait~0_combout ;


memory_control CC(
	.LessThan1(LessThan1),
	.always0(always0),
	.dhit(\CM|dhit~0_combout ),
	.iwait(\CC|iwait~0_combout ),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

caches CM(
	.dWEN_M(dWEN_M),
	.dREN_M(dREN_M),
	.dhit(\CM|dhit~0_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

datapath DP(
	.pc_out_3(pc_out_3),
	.pc_out_2(pc_out_2),
	.pc_out_5(pc_out_5),
	.pc_out_4(pc_out_4),
	.pc_out_7(pc_out_7),
	.pc_out_6(pc_out_6),
	.pc_out_9(pc_out_9),
	.pc_out_8(pc_out_8),
	.pc_out_11(pc_out_11),
	.pc_out_10(pc_out_10),
	.pc_out_13(pc_out_13),
	.pc_out_12(pc_out_12),
	.pc_out_15(pc_out_15),
	.pc_out_14(pc_out_14),
	.pc_out_17(pc_out_17),
	.pc_out_16(pc_out_16),
	.pc_out_19(pc_out_19),
	.pc_out_18(pc_out_18),
	.pc_out_21(pc_out_21),
	.pc_out_20(pc_out_20),
	.pc_out_23(pc_out_23),
	.pc_out_22(pc_out_22),
	.pc_out_25(pc_out_25),
	.pc_out_24(pc_out_24),
	.pc_out_27(pc_out_27),
	.pc_out_26(pc_out_26),
	.rdata2_M_0(rdata2_M_0),
	.rdata2_M_1(rdata2_M_1),
	.rdata2_M_2(rdata2_M_2),
	.rdata2_M_3(rdata2_M_3),
	.rdata2_M_4(rdata2_M_4),
	.rdata2_M_5(rdata2_M_5),
	.rdata2_M_6(rdata2_M_6),
	.rdata2_M_7(rdata2_M_7),
	.rdata2_M_8(rdata2_M_8),
	.rdata2_M_9(rdata2_M_9),
	.rdata2_M_10(rdata2_M_10),
	.rdata2_M_11(rdata2_M_11),
	.rdata2_M_12(rdata2_M_12),
	.rdata2_M_13(rdata2_M_13),
	.rdata2_M_14(rdata2_M_14),
	.rdata2_M_15(rdata2_M_15),
	.rdata2_M_16(rdata2_M_16),
	.rdata2_M_17(rdata2_M_17),
	.rdata2_M_18(rdata2_M_18),
	.rdata2_M_19(rdata2_M_19),
	.rdata2_M_20(rdata2_M_20),
	.rdata2_M_21(rdata2_M_21),
	.rdata2_M_22(rdata2_M_22),
	.rdata2_M_23(rdata2_M_23),
	.rdata2_M_24(rdata2_M_24),
	.rdata2_M_25(rdata2_M_25),
	.rdata2_M_26(rdata2_M_26),
	.rdata2_M_27(rdata2_M_27),
	.rdata2_M_28(rdata2_M_28),
	.rdata2_M_29(rdata2_M_29),
	.rdata2_M_30(rdata2_M_30),
	.rdata2_M_31(rdata2_M_31),
	.LessThan1(LessThan1),
	.porto_M_1(porto_M_1),
	.pc_out_1(pc_out_1),
	.dWEN_M1(dWEN_M),
	.dREN_M1(dREN_M),
	.porto_M_0(porto_M_0),
	.pc_out_0(pc_out_0),
	.porto_M_3(porto_M_3),
	.porto_M_2(porto_M_2),
	.porto_M_5(porto_M_5),
	.porto_M_4(porto_M_4),
	.porto_M_7(porto_M_7),
	.porto_M_6(porto_M_6),
	.porto_M_9(porto_M_9),
	.porto_M_8(porto_M_8),
	.porto_M_11(porto_M_11),
	.porto_M_10(porto_M_10),
	.porto_M_13(porto_M_13),
	.porto_M_12(porto_M_12),
	.porto_M_15(porto_M_15),
	.porto_M_14(porto_M_14),
	.porto_M_17(porto_M_17),
	.porto_M_16(porto_M_16),
	.porto_M_19(porto_M_19),
	.porto_M_18(porto_M_18),
	.porto_M_21(porto_M_21),
	.porto_M_20(porto_M_20),
	.porto_M_23(porto_M_23),
	.porto_M_22(porto_M_22),
	.porto_M_25(porto_M_25),
	.porto_M_24(porto_M_24),
	.porto_M_27(porto_M_27),
	.porto_M_26(porto_M_26),
	.porto_M_29(porto_M_29),
	.pc_out_29(pc_out_29),
	.porto_M_28(porto_M_28),
	.pc_out_28(pc_out_28),
	.porto_M_31(porto_M_31),
	.pc_out_31(pc_out_31),
	.porto_M_30(porto_M_30),
	.pc_out_30(pc_out_30),
	.always0(always0),
	.always1(always1),
	.\dpif.dmemload ({ramiframload_31,ramiframload_30,ramiframload_29,ramiframload_28,ramiframload_27,ramiframload_26,ramiframload_25,gnd,ramiframload_23,gnd,ramiframload_21,gnd,gnd,gnd,ramiframload_17,ramiframload_16,gnd,ramiframload_14,ramiframload_13,ramiframload_12,ramiframload_11,
ramiframload_10,gnd,ramiframload_8,gnd,ramiframload_6,gnd,gnd,gnd,ramiframload_2,ramiframload_1,ramiframload_0}),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_7(ramiframload_7),
	.ramiframload_9(ramiframload_9),
	.ramiframload_15(ramiframload_15),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_22(ramiframload_22),
	.ramiframload_24(ramiframload_24),
	.dhit(\CM|dhit~0_combout ),
	.iwait(\CC|iwait~0_combout ),
	.nRST(nRST),
	.nRST1(nRST1),
	.CLK(CLK),
	.halt_WB1(halt_WB),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module caches (
	dWEN_M,
	dREN_M,
	dhit,
	devpor,
	devclrn,
	devoe);
input 	dWEN_M;
input 	dREN_M;
output 	dhit;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X57_Y34_N28
cycloneive_lcell_comb \dhit~0 (
// Equation(s):
// dhit = (dREN_M1) # (dWEN_M1)

	.dataa(dREN_M),
	.datab(gnd),
	.datac(dWEN_M),
	.datad(gnd),
	.cin(gnd),
	.combout(dhit),
	.cout());
// synopsys translate_off
defparam \dhit~0 .lut_mask = 16'hFAFA;
defparam \dhit~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module datapath (
	pc_out_3,
	pc_out_2,
	pc_out_5,
	pc_out_4,
	pc_out_7,
	pc_out_6,
	pc_out_9,
	pc_out_8,
	pc_out_11,
	pc_out_10,
	pc_out_13,
	pc_out_12,
	pc_out_15,
	pc_out_14,
	pc_out_17,
	pc_out_16,
	pc_out_19,
	pc_out_18,
	pc_out_21,
	pc_out_20,
	pc_out_23,
	pc_out_22,
	pc_out_25,
	pc_out_24,
	pc_out_27,
	pc_out_26,
	rdata2_M_0,
	rdata2_M_1,
	rdata2_M_2,
	rdata2_M_3,
	rdata2_M_4,
	rdata2_M_5,
	rdata2_M_6,
	rdata2_M_7,
	rdata2_M_8,
	rdata2_M_9,
	rdata2_M_10,
	rdata2_M_11,
	rdata2_M_12,
	rdata2_M_13,
	rdata2_M_14,
	rdata2_M_15,
	rdata2_M_16,
	rdata2_M_17,
	rdata2_M_18,
	rdata2_M_19,
	rdata2_M_20,
	rdata2_M_21,
	rdata2_M_22,
	rdata2_M_23,
	rdata2_M_24,
	rdata2_M_25,
	rdata2_M_26,
	rdata2_M_27,
	rdata2_M_28,
	rdata2_M_29,
	rdata2_M_30,
	rdata2_M_31,
	LessThan1,
	porto_M_1,
	pc_out_1,
	dWEN_M1,
	dREN_M1,
	porto_M_0,
	pc_out_0,
	porto_M_3,
	porto_M_2,
	porto_M_5,
	porto_M_4,
	porto_M_7,
	porto_M_6,
	porto_M_9,
	porto_M_8,
	porto_M_11,
	porto_M_10,
	porto_M_13,
	porto_M_12,
	porto_M_15,
	porto_M_14,
	porto_M_17,
	porto_M_16,
	porto_M_19,
	porto_M_18,
	porto_M_21,
	porto_M_20,
	porto_M_23,
	porto_M_22,
	porto_M_25,
	porto_M_24,
	porto_M_27,
	porto_M_26,
	porto_M_29,
	pc_out_29,
	porto_M_28,
	pc_out_28,
	porto_M_31,
	pc_out_31,
	porto_M_30,
	pc_out_30,
	always0,
	always1,
	\dpif.dmemload ,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_7,
	ramiframload_9,
	ramiframload_15,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_22,
	ramiframload_24,
	dhit,
	iwait,
	nRST,
	nRST1,
	CLK,
	halt_WB1,
	devpor,
	devclrn,
	devoe);
output 	pc_out_3;
output 	pc_out_2;
output 	pc_out_5;
output 	pc_out_4;
output 	pc_out_7;
output 	pc_out_6;
output 	pc_out_9;
output 	pc_out_8;
output 	pc_out_11;
output 	pc_out_10;
output 	pc_out_13;
output 	pc_out_12;
output 	pc_out_15;
output 	pc_out_14;
output 	pc_out_17;
output 	pc_out_16;
output 	pc_out_19;
output 	pc_out_18;
output 	pc_out_21;
output 	pc_out_20;
output 	pc_out_23;
output 	pc_out_22;
output 	pc_out_25;
output 	pc_out_24;
output 	pc_out_27;
output 	pc_out_26;
output 	rdata2_M_0;
output 	rdata2_M_1;
output 	rdata2_M_2;
output 	rdata2_M_3;
output 	rdata2_M_4;
output 	rdata2_M_5;
output 	rdata2_M_6;
output 	rdata2_M_7;
output 	rdata2_M_8;
output 	rdata2_M_9;
output 	rdata2_M_10;
output 	rdata2_M_11;
output 	rdata2_M_12;
output 	rdata2_M_13;
output 	rdata2_M_14;
output 	rdata2_M_15;
output 	rdata2_M_16;
output 	rdata2_M_17;
output 	rdata2_M_18;
output 	rdata2_M_19;
output 	rdata2_M_20;
output 	rdata2_M_21;
output 	rdata2_M_22;
output 	rdata2_M_23;
output 	rdata2_M_24;
output 	rdata2_M_25;
output 	rdata2_M_26;
output 	rdata2_M_27;
output 	rdata2_M_28;
output 	rdata2_M_29;
output 	rdata2_M_30;
output 	rdata2_M_31;
input 	LessThan1;
output 	porto_M_1;
output 	pc_out_1;
output 	dWEN_M1;
output 	dREN_M1;
output 	porto_M_0;
output 	pc_out_0;
output 	porto_M_3;
output 	porto_M_2;
output 	porto_M_5;
output 	porto_M_4;
output 	porto_M_7;
output 	porto_M_6;
output 	porto_M_9;
output 	porto_M_8;
output 	porto_M_11;
output 	porto_M_10;
output 	porto_M_13;
output 	porto_M_12;
output 	porto_M_15;
output 	porto_M_14;
output 	porto_M_17;
output 	porto_M_16;
output 	porto_M_19;
output 	porto_M_18;
output 	porto_M_21;
output 	porto_M_20;
output 	porto_M_23;
output 	porto_M_22;
output 	porto_M_25;
output 	porto_M_24;
output 	porto_M_27;
output 	porto_M_26;
output 	porto_M_29;
output 	pc_out_29;
output 	porto_M_28;
output 	pc_out_28;
output 	porto_M_31;
output 	pc_out_31;
output 	porto_M_30;
output 	pc_out_30;
input 	always0;
input 	always1;
input 	[31:0] \dpif.dmemload ;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_7;
input 	ramiframload_9;
input 	ramiframload_15;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_22;
input 	ramiframload_24;
input 	dhit;
input 	iwait;
input 	nRST;
input 	nRST1;
input 	CLK;
output 	halt_WB1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \pc_when_branch[2]~1 ;
wire \pc_when_branch[2]~0_combout ;
wire \pc_when_branch[3]~3 ;
wire \pc_when_branch[3]~2_combout ;
wire \pc_plus_4[3]~2_combout ;
wire \pc_when_branch[4]~5 ;
wire \pc_when_branch[4]~4_combout ;
wire \pc_when_branch[5]~7 ;
wire \pc_when_branch[5]~6_combout ;
wire \pc_plus_4[4]~4_combout ;
wire \pc_plus_4[5]~6_combout ;
wire \pc_when_branch[6]~9 ;
wire \pc_when_branch[6]~8_combout ;
wire \pc_when_branch[7]~11 ;
wire \pc_when_branch[7]~10_combout ;
wire \pc_plus_4[6]~8_combout ;
wire \pc_when_branch[8]~13 ;
wire \pc_when_branch[8]~12_combout ;
wire \pc_when_branch[9]~15 ;
wire \pc_when_branch[9]~14_combout ;
wire \pc_plus_4[8]~12_combout ;
wire \pc_plus_4[9]~14_combout ;
wire \pc_when_branch[10]~17 ;
wire \pc_when_branch[10]~16_combout ;
wire \pc_when_branch[11]~19 ;
wire \pc_when_branch[11]~18_combout ;
wire \pc_plus_4[10]~16_combout ;
wire \pc_plus_4[11]~18_combout ;
wire \pc_when_branch[12]~21 ;
wire \pc_when_branch[12]~20_combout ;
wire \pc_when_branch[13]~23 ;
wire \pc_when_branch[13]~22_combout ;
wire \pc_plus_4[12]~20_combout ;
wire \pc_plus_4[13]~22_combout ;
wire \pc_when_branch[14]~25 ;
wire \pc_when_branch[14]~24_combout ;
wire \pc_when_branch[15]~27 ;
wire \pc_when_branch[15]~26_combout ;
wire \pc_plus_4[14]~24_combout ;
wire \pc_plus_4[15]~26_combout ;
wire \pc_when_branch[16]~29 ;
wire \pc_when_branch[16]~28_combout ;
wire \pc_when_branch[17]~31 ;
wire \pc_when_branch[17]~30_combout ;
wire \pc_plus_4[16]~28_combout ;
wire \pc_when_branch[18]~33 ;
wire \pc_when_branch[18]~32_combout ;
wire \pc_when_branch[19]~35 ;
wire \pc_when_branch[19]~34_combout ;
wire \pc_plus_4[18]~32_combout ;
wire \pc_when_branch[20]~37 ;
wire \pc_when_branch[20]~36_combout ;
wire \pc_when_branch[21]~39 ;
wire \pc_when_branch[21]~38_combout ;
wire \pc_plus_4[21]~38_combout ;
wire \pc_when_branch[22]~41 ;
wire \pc_when_branch[22]~40_combout ;
wire \pc_when_branch[23]~43 ;
wire \pc_when_branch[23]~42_combout ;
wire \pc_plus_4[22]~40_combout ;
wire \pc_when_branch[24]~45 ;
wire \pc_when_branch[24]~44_combout ;
wire \pc_when_branch[25]~47 ;
wire \pc_when_branch[25]~46_combout ;
wire \pc_plus_4[24]~44_combout ;
wire \pc_when_branch[26]~49 ;
wire \pc_when_branch[26]~48_combout ;
wire \pc_when_branch[27]~51 ;
wire \pc_when_branch[27]~50_combout ;
wire \pc_plus_4[26]~48_combout ;
wire \pc_plus_4[28]~52_combout ;
wire \pc_plus_4[29]~54_combout ;
wire \pc_when_branch[28]~53 ;
wire \pc_when_branch[28]~52_combout ;
wire \pc_when_branch[29]~55 ;
wire \pc_when_branch[29]~54_combout ;
wire \pc_plus_4[30]~57 ;
wire \pc_plus_4[31]~58_combout ;
wire \pc_when_branch[30]~57 ;
wire \pc_when_branch[30]~56_combout ;
wire \pc_when_branch[31]~58_combout ;
wire \Add2~1 ;
wire \Add2~0_combout ;
wire \Add2~3 ;
wire \Add2~2_combout ;
wire \Add2~5 ;
wire \Add2~4_combout ;
wire \Add2~7 ;
wire \Add2~6_combout ;
wire \Add2~9 ;
wire \Add2~8_combout ;
wire \Add2~11 ;
wire \Add2~10_combout ;
wire \Add2~13 ;
wire \Add2~12_combout ;
wire \Add2~15 ;
wire \Add2~14_combout ;
wire \Add2~17 ;
wire \Add2~16_combout ;
wire \Add2~19 ;
wire \Add2~18_combout ;
wire \Add2~21 ;
wire \Add2~20_combout ;
wire \Add2~23 ;
wire \Add2~22_combout ;
wire \Add2~25 ;
wire \Add2~24_combout ;
wire \Add2~27 ;
wire \Add2~26_combout ;
wire \Add2~29 ;
wire \Add2~28_combout ;
wire \Add2~31 ;
wire \Add2~30_combout ;
wire \Add2~33 ;
wire \Add2~32_combout ;
wire \Add2~35 ;
wire \Add2~34_combout ;
wire \Add2~37 ;
wire \Add2~36_combout ;
wire \Add2~39 ;
wire \Add2~38_combout ;
wire \Add2~41 ;
wire \Add2~40_combout ;
wire \Add2~43 ;
wire \Add2~42_combout ;
wire \Add2~45 ;
wire \Add2~44_combout ;
wire \Add2~47 ;
wire \Add2~46_combout ;
wire \Add2~49 ;
wire \Add2~48_combout ;
wire \Add2~51 ;
wire \Add2~50_combout ;
wire \Add2~53 ;
wire \Add2~52_combout ;
wire \Add2~55 ;
wire \Add2~54_combout ;
wire \Add2~57 ;
wire \Add2~56_combout ;
wire \Add2~58_combout ;
wire \rdata1_M[1]~31_combout ;
wire \rdata1_M[0]~30_combout ;
wire \rdata1_M[3]~0_combout ;
wire \rdata1_M[2]~1_combout ;
wire \rdata1_M[5]~3_combout ;
wire \rdata1_M[4]~2_combout ;
wire \rdata1_M[7]~5_combout ;
wire \rdata1_M[6]~4_combout ;
wire \rdata1_M[9]~7_combout ;
wire \rdata1_M[8]~6_combout ;
wire \rdata1_M[11]~9_combout ;
wire \rdata1_M[10]~8_combout ;
wire \rdata1_M[13]~11_combout ;
wire \rdata1_M[12]~10_combout ;
wire \rdata1_M[15]~13_combout ;
wire \rdata1_M[14]~12_combout ;
wire \rdata1_M[17]~15_combout ;
wire \rdata1_M[16]~14_combout ;
wire \rdata1_M[19]~17_combout ;
wire \rdata1_M[18]~16_combout ;
wire \rdata1_M[21]~19_combout ;
wire \rdata1_M[20]~18_combout ;
wire \rdata1_M[23]~21_combout ;
wire \rdata1_M[22]~20_combout ;
wire \rdata1_M[25]~23_combout ;
wire \rdata1_M[24]~22_combout ;
wire \rdata1_M[27]~25_combout ;
wire \rdata1_M[26]~24_combout ;
wire \rdata1_M[29]~27_combout ;
wire \rdata1_M[28]~26_combout ;
wire \rdata1_M[31]~29_combout ;
wire \rdata1_M[30]~28_combout ;
wire \bne_M~q ;
wire \jr_M~q ;
wire \Equal4~0_combout ;
wire \Equal4~1_combout ;
wire \FORWARDING_UNIT|Equal0~2_combout ;
wire \FORWARDING_UNIT|fuif.forward_A[0]~2_combout ;
wire \FORWARDING_UNIT|fuif.forward_A[1]~5_combout ;
wire \FORWARDING_UNIT|fuif.bubble_lw_f~2_combout ;
wire \FORWARDING_UNIT|forward_B~0_combout ;
wire \beq_EX~q ;
wire \bne_EX~q ;
wire \FORWARDING_UNIT|forward_B~1_combout ;
wire \FORWARDING_UNIT|Equal5~1_combout ;
wire \ALUSrc_EX~q ;
wire \FORWARDING_UNIT|fuif.forward_B[1]~3_combout ;
wire \FORWARDING_UNIT|fuif.forward_B[1]~4_combout ;
wire \portB~15_combout ;
wire \portB~16_combout ;
wire \portB~17_combout ;
wire \portB~27_combout ;
wire \portB~28_combout ;
wire \portB~29_combout ;
wire \sw_forwarding_output~5_combout ;
wire \portB~33_combout ;
wire \portB~34_combout ;
wire \portB~35_combout ;
wire \portB~36_combout ;
wire \portB~37_combout ;
wire \portB~38_combout ;
wire \portB~39_combout ;
wire \portB~40_combout ;
wire \portB~41_combout ;
wire \portB~42_combout ;
wire \sw_forwarding_output~9_combout ;
wire \portB~43_combout ;
wire \portB~44_combout ;
wire \portB~48_combout ;
wire \portB~49_combout ;
wire \portB~50_combout ;
wire \portB~57_combout ;
wire \portB~58_combout ;
wire \portB~59_combout ;
wire \portB~60_combout ;
wire \sw_forwarding_output~17_combout ;
wire \portB~67_combout ;
wire \portB~68_combout ;
wire \portB~69_combout ;
wire \portB~70_combout ;
wire \portB~74_combout ;
wire \portB~75_combout ;
wire \portB~76_combout ;
wire \portB~77_combout ;
wire \portB~78_combout ;
wire \portB~79_combout ;
wire \portB~80_combout ;
wire \portB~81_combout ;
wire \portB~82_combout ;
wire \sw_forwarding_output~25_combout ;
wire \portB~85_combout ;
wire \portB~86_combout ;
wire \portB~87_combout ;
wire \FORWARDING_UNIT|Equal3~0_combout ;
wire \FORWARDING_UNIT|fuif.forward_A[0]~6_combout ;
wire \portA~8_combout ;
wire \FORWARDING_UNIT|Equal3~1_combout ;
wire \FORWARDING_UNIT|fuif.forward_A[1]~7_combout ;
wire \portA~9_combout ;
wire \portA~10_combout ;
wire \portA~11_combout ;
wire \portA~12_combout ;
wire \portB~89_combout ;
wire \portB~90_combout ;
wire \portB~91_combout ;
wire \portB~92_combout ;
wire \portB~94_combout ;
wire \portB~95_combout ;
wire \portB~96_combout ;
wire \portB~97_combout ;
wire \wdat_WB[4]~62_combout ;
wire \portA~13_combout ;
wire \portA~14_combout ;
wire \portA~15_combout ;
wire \portA~16_combout ;
wire \portA~17_combout ;
wire \portA~18_combout ;
wire \portA~19_combout ;
wire \portA~20_combout ;
wire \portA~21_combout ;
wire \portA~22_combout ;
wire \portA~23_combout ;
wire \portB~101_combout ;
wire \portB~102_combout ;
wire \portB~103_combout ;
wire \portA~24_combout ;
wire \portA~25_combout ;
wire \portA~26_combout ;
wire \portA~27_combout ;
wire \portA~28_combout ;
wire \portA~29_combout ;
wire \portA~30_combout ;
wire \portA~31_combout ;
wire \portA~32_combout ;
wire \portA~33_combout ;
wire \portA~34_combout ;
wire \portA~35_combout ;
wire \portA~36_combout ;
wire \portA~37_combout ;
wire \portA~38_combout ;
wire \portA~39_combout ;
wire \portA~40_combout ;
wire \portA~41_combout ;
wire \portA~42_combout ;
wire \portA~43_combout ;
wire \portA~44_combout ;
wire \portA~45_combout ;
wire \portA~46_combout ;
wire \portA~47_combout ;
wire \portA~48_combout ;
wire \portA~49_combout ;
wire \portA~50_combout ;
wire \portA~51_combout ;
wire \portA~52_combout ;
wire \portA~53_combout ;
wire \portA~54_combout ;
wire \portA~55_combout ;
wire \portA~56_combout ;
wire \portA~57_combout ;
wire \portA~58_combout ;
wire \portA~59_combout ;
wire \portA~60_combout ;
wire \portA~61_combout ;
wire \portA~62_combout ;
wire \portA~63_combout ;
wire \portA~64_combout ;
wire \portA~65_combout ;
wire \portA~66_combout ;
wire \portA~67_combout ;
wire \ALU|Selector0~5_combout ;
wire \ALU|Selector30~8_combout ;
wire \pc_next[1]~0_combout ;
wire \pc_next[1]~1_combout ;
wire \pc_next[1]~2_combout ;
wire \btbframes.frameblocks[2].valid~q ;
wire \btbframes.frameblocks[1].valid~q ;
wire \btbframes.frameblocks[0].valid~q ;
wire \btbframes.frameblocks[3].valid~q ;
wire \BTB|predicted~18_combout ;
wire \pc_next~3_combout ;
wire \pc_next[1]~4_combout ;
wire \CONTROL_UNIT|Decoder1~0_combout ;
wire \CONTROL_UNIT|Decoder1~1_combout ;
wire \portB~108_combout ;
wire \portB~109_combout ;
wire \ALU|Selector31~4_combout ;
wire \ALU|Selector31~5_combout ;
wire \ALU|Selector31~8_combout ;
wire \pc_next[0]~5_combout ;
wire \pc_next[0]~6_combout ;
wire \pc_next[0]~7_combout ;
wire \pc_next[0]~8_combout ;
wire \ALU|Selector28~10_combout ;
wire \pc_next[3]~9_combout ;
wire \pc_next[3]~10_combout ;
wire \pc_next[3]~11_combout ;
wire \pc_next[3]~12_combout ;
wire \comb~2_combout ;
wire \ALU|Selector29~10_combout ;
wire \pc_next[2]~13_combout ;
wire \pc_next[2]~14_combout ;
wire \pc_next[2]~15_combout ;
wire \pc_next[2]~16_combout ;
wire \ALU|Selector26~6_combout ;
wire \pc_next[5]~17_combout ;
wire \pc_next[5]~18_combout ;
wire \pc_next[5]~19_combout ;
wire \pc_next[5]~20_combout ;
wire \ALU|Selector27~0_combout ;
wire \ALU|Selector27~3_combout ;
wire \ALU|Selector27~6_combout ;
wire \ALU|Selector27~7_combout ;
wire \pc_next[4]~21_combout ;
wire \pc_next[4]~22_combout ;
wire \pc_next[4]~23_combout ;
wire \pc_next[4]~24_combout ;
wire \ALU|Selector24~8_combout ;
wire \pc_next[7]~25_combout ;
wire \pc_next[7]~26_combout ;
wire \pc_next[7]~27_combout ;
wire \pc_next[7]~28_combout ;
wire \ALU|Selector25~7_combout ;
wire \pc_next[6]~29_combout ;
wire \pc_next[6]~30_combout ;
wire \pc_next[6]~31_combout ;
wire \pc_next[6]~32_combout ;
wire \ALU|Selector22~8_combout ;
wire \pc_next[9]~33_combout ;
wire \pc_next[9]~34_combout ;
wire \pc_next[9]~35_combout ;
wire \pc_next[9]~36_combout ;
wire \ALU|Selector16~3_combout ;
wire \ALU|Selector23~8_combout ;
wire \pc_next[8]~37_combout ;
wire \pc_next[8]~38_combout ;
wire \pc_next[8]~39_combout ;
wire \pc_next[8]~40_combout ;
wire \ALU|Selector20~8_combout ;
wire \pc_next[11]~41_combout ;
wire \pc_next[11]~42_combout ;
wire \pc_next[11]~43_combout ;
wire \pc_next[11]~44_combout ;
wire \ALU|Selector21~7_combout ;
wire \pc_next[10]~45_combout ;
wire \pc_next[10]~46_combout ;
wire \pc_next[10]~47_combout ;
wire \pc_next[10]~48_combout ;
wire \ALU|Selector18~7_combout ;
wire \pc_next[13]~49_combout ;
wire \pc_next[13]~50_combout ;
wire \pc_next[13]~51_combout ;
wire \pc_next[13]~52_combout ;
wire \ALU|Selector19~6_combout ;
wire \ALU|ShiftLeft0~57_combout ;
wire \pc_next[12]~53_combout ;
wire \pc_next[12]~54_combout ;
wire \pc_next[12]~55_combout ;
wire \pc_next[12]~56_combout ;
wire \ALU|Selector16~11_combout ;
wire \pc_next[15]~57_combout ;
wire \pc_next[15]~58_combout ;
wire \pc_next[15]~59_combout ;
wire \pc_next[15]~60_combout ;
wire \ALU|Selector17~8_combout ;
wire \pc_next[14]~61_combout ;
wire \pc_next[14]~62_combout ;
wire \pc_next[14]~63_combout ;
wire \pc_next[14]~64_combout ;
wire \ALU|Selector12~10_combout ;
wire \ALU|Selector14~7_combout ;
wire \pc_next[17]~65_combout ;
wire \pc_next[17]~66_combout ;
wire \pc_next[17]~67_combout ;
wire \pc_next[17]~68_combout ;
wire \ALU|Selector15~11_combout ;
wire \pc_next[16]~69_combout ;
wire \pc_next[16]~70_combout ;
wire \pc_next[16]~71_combout ;
wire \pc_next[16]~72_combout ;
wire \ALU|Selector12~18_combout ;
wire \pc_next[19]~73_combout ;
wire \pc_next[19]~74_combout ;
wire \pc_next[19]~75_combout ;
wire \pc_next[19]~76_combout ;
wire \ALU|Selector13~8_combout ;
wire \pc_next[18]~77_combout ;
wire \pc_next[18]~78_combout ;
wire \pc_next[18]~79_combout ;
wire \pc_next[18]~80_combout ;
wire \ALU|Selector10~8_combout ;
wire \pc_next[21]~81_combout ;
wire \pc_next[21]~82_combout ;
wire \pc_next[21]~83_combout ;
wire \pc_next[21]~84_combout ;
wire \ALU|Selector11~8_combout ;
wire \pc_next[20]~85_combout ;
wire \pc_next[20]~86_combout ;
wire \pc_next[20]~87_combout ;
wire \pc_next[20]~88_combout ;
wire \ALU|Selector8~7_combout ;
wire \pc_next[23]~89_combout ;
wire \pc_next[23]~90_combout ;
wire \pc_next[23]~91_combout ;
wire \pc_next[23]~92_combout ;
wire \ALU|Selector9~8_combout ;
wire \pc_next[22]~93_combout ;
wire \pc_next[22]~94_combout ;
wire \pc_next[22]~95_combout ;
wire \pc_next[22]~96_combout ;
wire \ALU|Selector6~0_combout ;
wire \ALU|Selector6~5_combout ;
wire \ALU|Selector6~7_combout ;
wire \pc_next[25]~97_combout ;
wire \pc_next[25]~98_combout ;
wire \pc_next[25]~99_combout ;
wire \pc_next[25]~100_combout ;
wire \ALU|Selector7~7_combout ;
wire \pc_next[24]~101_combout ;
wire \pc_next[24]~102_combout ;
wire \pc_next[24]~103_combout ;
wire \pc_next[24]~104_combout ;
wire \ALU|Selector4~12_combout ;
wire \pc_next[27]~105_combout ;
wire \pc_next[27]~106_combout ;
wire \pc_next[27]~107_combout ;
wire \pc_next[27]~108_combout ;
wire \ALU|Selector5~7_combout ;
wire \pc_next[26]~109_combout ;
wire \pc_next[26]~110_combout ;
wire \pc_next[26]~111_combout ;
wire \pc_next[26]~112_combout ;
wire \ALU|Selector2~11_combout ;
wire \pc_next[29]~113_combout ;
wire \pc_next[29]~114_combout ;
wire \PROGRAM_COUNTER|pc_out[29]~29_combout ;
wire \PROGRAM_COUNTER|pc_out[29]~30_combout ;
wire \pc_next[29]~115_combout ;
wire \pc_next[29]~116_combout ;
wire \pc_next[29]~117_combout ;
wire \ALU|Selector3~9_combout ;
wire \pc_next[28]~118_combout ;
wire \pc_next[28]~119_combout ;
wire \pc_next[28]~120_combout ;
wire \pc_next[28]~121_combout ;
wire \pc_next[28]~122_combout ;
wire \ALU|Selector0~27_combout ;
wire \pc_next[31]~123_combout ;
wire \pc_next[31]~124_combout ;
wire \pc_next[31]~125_combout ;
wire \pc_next[31]~126_combout ;
wire \pc_next[31]~127_combout ;
wire \ALU|Selector1~9_combout ;
wire \pc_next[30]~128_combout ;
wire \pc_next[30]~129_combout ;
wire \pc_next[30]~130_combout ;
wire \pc_next[30]~131_combout ;
wire \pc_next[30]~132_combout ;
wire \cu_halt_EX~q ;
wire \jal_EX~q ;
wire \predicted_EX~q ;
wire \bne_M~0_combout ;
wire \ALU|Selector6~8_combout ;
wire \ALU|Selector6~9_combout ;
wire \zero_M~5_combout ;
wire \ALU|Selector31~9_combout ;
wire \jr_EX~q ;
wire \jr_M~0_combout ;
wire \op_EX~0_combout ;
wire \op_EX~1_combout ;
wire \op_EX~2_combout ;
wire \op_EX~3_combout ;
wire \op_EX~4_combout ;
wire \op_EX~5_combout ;
wire \instruction_EX~0_combout ;
wire \instruction_EX~1_combout ;
wire \RegDst_EX~q ;
wire \wsel_M~1_combout ;
wire \wsel_M~2_combout ;
wire \wsel_M~3_combout ;
wire \wsel_M~4_combout ;
wire \instruction_EX~2_combout ;
wire \instruction_EX~3_combout ;
wire \wsel_M~5_combout ;
wire \wsel_M~6_combout ;
wire \wsel_M~7_combout ;
wire \wsel_M~8_combout ;
wire \instruction_EX~4_combout ;
wire \wsel_M~9_combout ;
wire \wsel_M~10_combout ;
wire \instruction_EX~5_combout ;
wire \instruction_EX~7_combout ;
wire \instruction_EX~8_combout ;
wire \instruction_EX~9_combout ;
wire \CONTROL_UNIT|Equal3~1_combout ;
wire \CONTROL_UNIT|Equal3~2_combout ;
wire \CONTROL_UNIT|WideOr2~0_combout ;
wire \ALUOp_EX~0_combout ;
wire \ALUOp_EX~1_combout ;
wire \CONTROL_UNIT|WideOr7~0_combout ;
wire \ALUOp_EX~2_combout ;
wire \ALUOp_EX~3_combout ;
wire \CONTROL_UNIT|WideOr6~0_combout ;
wire \ALUOp_EX~4_combout ;
wire \ALUOp_EX~5_combout ;
wire \CONTROL_UNIT|WideOr1~0_combout ;
wire \ALUOp_EX~6_combout ;
wire \ALUOp_EX~7_combout ;
wire \ALUOp_EX~8_combout ;
wire \ALUOp_EX~9_combout ;
wire \CONTROL_UNIT|WideOr5~0_combout ;
wire \ALUOp_EX~10_combout ;
wire \ALUOp_EX~11_combout ;
wire \ALUOp_EX~12_combout ;
wire \ALUOp_EX~13_combout ;
wire \ExtOp_EX~0_combout ;
wire \CONTROL_UNIT|WideOr8~0_combout ;
wire \RegWrite_EX~q ;
wire \beq_EX~0_combout ;
wire \bne_EX~0_combout ;
wire \CONTROL_UNIT|WideOr4~0_combout ;
wire \ALUSrc_EX~1_combout ;
wire \REGISTER_FILE|Mux32~9_combout ;
wire \REGISTER_FILE|Mux32~19_combout ;
wire \lui_EX~q ;
wire \REGISTER_FILE|Mux33~9_combout ;
wire \REGISTER_FILE|Mux33~19_combout ;
wire \REGISTER_FILE|Mux34~9_combout ;
wire \REGISTER_FILE|Mux34~19_combout ;
wire \REGISTER_FILE|Mux35~9_combout ;
wire \REGISTER_FILE|Mux35~19_combout ;
wire \REGISTER_FILE|Mux36~9_combout ;
wire \REGISTER_FILE|Mux36~19_combout ;
wire \rdata2_EX~8_combout ;
wire \rdata2_EX~9_combout ;
wire \REGISTER_FILE|Mux37~9_combout ;
wire \REGISTER_FILE|Mux37~19_combout ;
wire \REGISTER_FILE|Mux38~9_combout ;
wire \REGISTER_FILE|Mux38~19_combout ;
wire \rdata2_EX~12_combout ;
wire \rdata2_EX~13_combout ;
wire \REGISTER_FILE|Mux39~9_combout ;
wire \REGISTER_FILE|Mux39~19_combout ;
wire \REGISTER_FILE|Mux40~9_combout ;
wire \REGISTER_FILE|Mux40~19_combout ;
wire \REGISTER_FILE|Mux41~9_combout ;
wire \REGISTER_FILE|Mux41~19_combout ;
wire \REGISTER_FILE|Mux42~9_combout ;
wire \REGISTER_FILE|Mux42~19_combout ;
wire \REGISTER_FILE|Mux43~9_combout ;
wire \REGISTER_FILE|Mux43~19_combout ;
wire \rdata2_EX~22_combout ;
wire \rdata2_EX~23_combout ;
wire \REGISTER_FILE|Mux44~9_combout ;
wire \REGISTER_FILE|Mux44~19_combout ;
wire \REGISTER_FILE|Mux45~9_combout ;
wire \REGISTER_FILE|Mux45~19_combout ;
wire \REGISTER_FILE|Mux46~9_combout ;
wire \REGISTER_FILE|Mux46~19_combout ;
wire \REGISTER_FILE|Mux47~9_combout ;
wire \REGISTER_FILE|Mux47~19_combout ;
wire \REGISTER_FILE|Mux48~9_combout ;
wire \REGISTER_FILE|Mux48~19_combout ;
wire \REGISTER_FILE|Mux49~9_combout ;
wire \REGISTER_FILE|Mux49~19_combout ;
wire \REGISTER_FILE|Mux50~9_combout ;
wire \REGISTER_FILE|Mux50~19_combout ;
wire \rdata2_EX~36_combout ;
wire \rdata2_EX~37_combout ;
wire \REGISTER_FILE|Mux51~9_combout ;
wire \REGISTER_FILE|Mux51~19_combout ;
wire \REGISTER_FILE|Mux54~9_combout ;
wire \REGISTER_FILE|Mux54~19_combout ;
wire \REGISTER_FILE|Mux55~9_combout ;
wire \REGISTER_FILE|Mux55~19_combout ;
wire \rdata2_EX~42_combout ;
wire \rdata2_EX~43_combout ;
wire \imm_EX~6_combout ;
wire \REGISTER_FILE|Mux52~9_combout ;
wire \REGISTER_FILE|Mux52~19_combout ;
wire \rdata2_EX~44_combout ;
wire \rdata2_EX~45_combout ;
wire \REGISTER_FILE|Mux53~9_combout ;
wire \REGISTER_FILE|Mux53~19_combout ;
wire \rdata2_EX~46_combout ;
wire \rdata2_EX~47_combout ;
wire \REGISTER_FILE|Mux56~9_combout ;
wire \REGISTER_FILE|Mux56~19_combout ;
wire \rdata2_EX~48_combout ;
wire \rdata2_EX~49_combout ;
wire \REGISTER_FILE|Mux57~9_combout ;
wire \REGISTER_FILE|Mux57~19_combout ;
wire \REGISTER_FILE|Mux58~9_combout ;
wire \REGISTER_FILE|Mux58~19_combout ;
wire \rdata2_EX~52_combout ;
wire \rdata2_EX~53_combout ;
wire \REGISTER_FILE|Mux29~9_combout ;
wire \REGISTER_FILE|Mux29~19_combout ;
wire \rdata1_EX~2_combout ;
wire \rdata1_EX~3_combout ;
wire \REGISTER_FILE|Mux30~9_combout ;
wire \REGISTER_FILE|Mux30~19_combout ;
wire \rdata1_EX~4_combout ;
wire \rdata1_EX~5_combout ;
wire \REGISTER_FILE|Mux63~9_combout ;
wire \REGISTER_FILE|Mux63~19_combout ;
wire \rdata2_EX~54_combout ;
wire \rdata2_EX~55_combout ;
wire \REGISTER_FILE|Mux62~9_combout ;
wire \REGISTER_FILE|Mux62~19_combout ;
wire \rdata2_EX~56_combout ;
wire \rdata2_EX~57_combout ;
wire \REGISTER_FILE|Mux27~9_combout ;
wire \REGISTER_FILE|Mux27~19_combout ;
wire \rdata1_EX~6_combout ;
wire \rdata1_EX~7_combout ;
wire \REGISTER_FILE|Mux28~9_combout ;
wire \REGISTER_FILE|Mux28~19_combout ;
wire \rdata1_EX~8_combout ;
wire \rdata1_EX~9_combout ;
wire \REGISTER_FILE|Mux61~9_combout ;
wire \REGISTER_FILE|Mux61~19_combout ;
wire \REGISTER_FILE|Mux23~9_combout ;
wire \REGISTER_FILE|Mux23~19_combout ;
wire \rdata1_EX~10_combout ;
wire \rdata1_EX~11_combout ;
wire \REGISTER_FILE|Mux24~9_combout ;
wire \REGISTER_FILE|Mux24~19_combout ;
wire \rdata1_EX~12_combout ;
wire \rdata1_EX~13_combout ;
wire \REGISTER_FILE|Mux25~9_combout ;
wire \REGISTER_FILE|Mux25~19_combout ;
wire \rdata1_EX~14_combout ;
wire \rdata1_EX~15_combout ;
wire \REGISTER_FILE|Mux26~9_combout ;
wire \REGISTER_FILE|Mux26~19_combout ;
wire \rdata1_EX~16_combout ;
wire \rdata1_EX~17_combout ;
wire \REGISTER_FILE|Mux60~9_combout ;
wire \REGISTER_FILE|Mux60~19_combout ;
wire \rdata2_EX~60_combout ;
wire \rdata2_EX~61_combout ;
wire \REGISTER_FILE|Mux15~9_combout ;
wire \REGISTER_FILE|Mux15~19_combout ;
wire \rdata1_EX~18_combout ;
wire \rdata1_EX~19_combout ;
wire \REGISTER_FILE|Mux16~9_combout ;
wire \REGISTER_FILE|Mux16~19_combout ;
wire \rdata1_EX~20_combout ;
wire \rdata1_EX~21_combout ;
wire \REGISTER_FILE|Mux17~9_combout ;
wire \REGISTER_FILE|Mux17~19_combout ;
wire \rdata1_EX~22_combout ;
wire \rdata1_EX~23_combout ;
wire \REGISTER_FILE|Mux18~9_combout ;
wire \REGISTER_FILE|Mux18~19_combout ;
wire \rdata1_EX~24_combout ;
wire \rdata1_EX~25_combout ;
wire \REGISTER_FILE|Mux19~9_combout ;
wire \REGISTER_FILE|Mux19~19_combout ;
wire \rdata1_EX~26_combout ;
wire \rdata1_EX~27_combout ;
wire \REGISTER_FILE|Mux20~9_combout ;
wire \REGISTER_FILE|Mux20~19_combout ;
wire \rdata1_EX~28_combout ;
wire \rdata1_EX~29_combout ;
wire \REGISTER_FILE|Mux21~9_combout ;
wire \REGISTER_FILE|Mux21~19_combout ;
wire \rdata1_EX~30_combout ;
wire \rdata1_EX~31_combout ;
wire \REGISTER_FILE|Mux22~9_combout ;
wire \REGISTER_FILE|Mux22~19_combout ;
wire \rdata1_EX~32_combout ;
wire \rdata1_EX~33_combout ;
wire \REGISTER_FILE|Mux59~9_combout ;
wire \REGISTER_FILE|Mux59~19_combout ;
wire \REGISTER_FILE|Mux0~9_combout ;
wire \REGISTER_FILE|Mux0~19_combout ;
wire \rdata1_EX~34_combout ;
wire \rdata1_EX~35_combout ;
wire \REGISTER_FILE|Mux2~9_combout ;
wire \REGISTER_FILE|Mux2~19_combout ;
wire \rdata1_EX~36_combout ;
wire \rdata1_EX~37_combout ;
wire \REGISTER_FILE|Mux1~9_combout ;
wire \REGISTER_FILE|Mux1~19_combout ;
wire \rdata1_EX~38_combout ;
wire \rdata1_EX~39_combout ;
wire \REGISTER_FILE|Mux3~9_combout ;
wire \REGISTER_FILE|Mux3~19_combout ;
wire \rdata1_EX~40_combout ;
wire \rdata1_EX~41_combout ;
wire \REGISTER_FILE|Mux4~9_combout ;
wire \REGISTER_FILE|Mux4~19_combout ;
wire \rdata1_EX~42_combout ;
wire \rdata1_EX~43_combout ;
wire \REGISTER_FILE|Mux5~9_combout ;
wire \REGISTER_FILE|Mux5~19_combout ;
wire \rdata1_EX~44_combout ;
wire \rdata1_EX~45_combout ;
wire \REGISTER_FILE|Mux6~9_combout ;
wire \REGISTER_FILE|Mux6~19_combout ;
wire \rdata1_EX~46_combout ;
wire \rdata1_EX~47_combout ;
wire \REGISTER_FILE|Mux7~9_combout ;
wire \REGISTER_FILE|Mux7~19_combout ;
wire \rdata1_EX~48_combout ;
wire \rdata1_EX~49_combout ;
wire \REGISTER_FILE|Mux8~9_combout ;
wire \REGISTER_FILE|Mux8~19_combout ;
wire \rdata1_EX~50_combout ;
wire \rdata1_EX~51_combout ;
wire \REGISTER_FILE|Mux9~9_combout ;
wire \REGISTER_FILE|Mux9~19_combout ;
wire \rdata1_EX~52_combout ;
wire \rdata1_EX~53_combout ;
wire \REGISTER_FILE|Mux10~9_combout ;
wire \REGISTER_FILE|Mux10~19_combout ;
wire \rdata1_EX~54_combout ;
wire \rdata1_EX~55_combout ;
wire \REGISTER_FILE|Mux11~9_combout ;
wire \REGISTER_FILE|Mux11~19_combout ;
wire \rdata1_EX~56_combout ;
wire \rdata1_EX~57_combout ;
wire \REGISTER_FILE|Mux12~9_combout ;
wire \REGISTER_FILE|Mux12~19_combout ;
wire \rdata1_EX~58_combout ;
wire \rdata1_EX~59_combout ;
wire \REGISTER_FILE|Mux13~9_combout ;
wire \REGISTER_FILE|Mux13~19_combout ;
wire \rdata1_EX~60_combout ;
wire \rdata1_EX~61_combout ;
wire \REGISTER_FILE|Mux14~9_combout ;
wire \REGISTER_FILE|Mux14~19_combout ;
wire \rdata1_EX~62_combout ;
wire \rdata1_EX~63_combout ;
wire \REGISTER_FILE|Mux31~9_combout ;
wire \REGISTER_FILE|Mux31~19_combout ;
wire \Decoder0~0_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \does_exist~0_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \does_exist~1_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \does_exist~2_combout ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \does_exist~3_combout ;
wire \does_exist~4_combout ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \does_exist~5_combout ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \does_exist~6_combout ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \does_exist~7_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \does_exist~8_combout ;
wire \always3~2_combout ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \does_exist~9_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \does_exist~10_combout ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \does_exist~11_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \does_exist~12_combout ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \does_exist~13_combout ;
wire \does_exist~14_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \does_exist~15_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \does_exist~16_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \does_exist~17_combout ;
wire \does_exist~18_combout ;
wire \btbframes.frameblocks[2].tag[27]~2_combout ;
wire \Decoder0~1_combout ;
wire \btbframes.frameblocks[1].tag[27]~2_combout ;
wire \btbframes.frameblocks[0].tag[27]~2_combout ;
wire \Decoder0~2_combout ;
wire \btbframes.frameblocks[3].tag[27]~2_combout ;
wire \rdata1_M~32_combout ;
wire \rdata1_M~33_combout ;
wire \btbframes.frameblocks[0].valid~0_combout ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \btbframes~0_combout ;
wire \btbframes~1_combout ;
wire \btbframes.frameblocks[2].curr_state[0]~0_combout ;
wire \btbframes.frameblocks[2].curr_state[0]~1_combout ;
wire \btbframes.frameblocks[1].curr_state[1]~0_combout ;
wire \btbframes.frameblocks[1].curr_state[1]~1_combout ;
wire \btbframes.frameblocks[2].curr_state[1]~2_combout ;
wire \btbframes.frameblocks[1].curr_state[1]~2_combout ;
wire \btbframes.frameblocks[2].curr_state[1]~3_combout ;
wire \btbframes.frameblocks[0].curr_state[1]~0_combout ;
wire \btbframes.frameblocks[0].curr_state[1]~1_combout ;
wire \btbframes.frameblocks[0].curr_state[1]~2_combout ;
wire \btbframes.frameblocks[3].curr_state[1]~0_combout ;
wire \pc_plus_4_M~17_combout ;
wire \pc_plus_4_M~19_combout ;
wire \instruction_M~0_combout ;
wire \instruction_M~1_combout ;
wire \pc_plus_4_M~20_combout ;
wire \instruction_M~2_combout ;
wire \instruction_M~3_combout ;
wire \instruction_M~4_combout ;
wire \instruction_M~5_combout ;
wire \instruction_M~6_combout ;
wire \instruction_M~7_combout ;
wire \instruction_M~8_combout ;
wire \instruction_M~9_combout ;
wire \pc_plus_4_M~29_combout ;
wire \sw_forwarding_output~29_combout ;
wire \sw_forwarding_output~31_combout ;
wire \cu_halt_EX~0_combout ;
wire \predicted_D~q ;
wire \predicted_EX~0_combout ;
wire \CONTROL_UNIT|Decoder0~1_combout ;
wire \jr_EX~0_combout ;
wire \op_D~0_combout ;
wire \op_D~1_combout ;
wire \op_D~2_combout ;
wire \op_D~3_combout ;
wire \op_D~4_combout ;
wire \op_D~5_combout ;
wire \op_D~6_combout ;
wire \op_D~7_combout ;
wire \op_D~8_combout ;
wire \op_D~9_combout ;
wire \op_D~10_combout ;
wire \op_D~11_combout ;
wire \RegDst_EX~0_combout ;
wire \RegWrite_EX~0_combout ;
wire \RegWrite_EX~1_combout ;
wire \RegWrite_EX~2_combout ;
wire \RegWrite_EX~3_combout ;
wire \lui_EX~1_combout ;
wire \pc_plus_4_EX~0_combout ;
wire \btbframes~2_combout ;
wire \btbframes.frameblocks[3].curr_state[0]~1_combout ;
wire \btbframes.frameblocks[3].curr_state[0]~2_combout ;
wire \btbframes.frameblocks[2].curr_state[0]~4_combout ;
wire \btbframes.frameblocks[1].curr_state[0]~3_combout ;
wire \btbframes.frameblocks[0].curr_state[0]~3_combout ;
wire \btbframes.frameblocks[3].curr_state[0]~3_combout ;
wire \pc_plus_4_EX~9_combout ;
wire \pc_plus_4_EX~13_combout ;
wire \pc_plus_4_EX~14_combout ;
wire \pc_plus_4_EX~15_combout ;
wire \pc_plus_4_EX~17_combout ;
wire \pc_plus_4_EX~19_combout ;
wire \pc_plus_4_EX~20_combout ;
wire \pc_plus_4_EX~23_combout ;
wire \pc_plus_4_EX~28_combout ;
wire \pc_plus_4_EX~29_combout ;
wire \predicted_D~0_combout ;
wire \pc_plus_4_D~0_combout ;
wire \pc_plus_4_D~2_combout ;
wire \pc_plus_4_D~4_combout ;
wire \pc_plus_4_D~5_combout ;
wire \pc_plus_4_D~7_combout ;
wire \pc_plus_4_D~8_combout ;
wire \pc_plus_4_D~9_combout ;
wire \pc_plus_4_D~10_combout ;
wire \pc_plus_4_D~11_combout ;
wire \pc_plus_4_D~12_combout ;
wire \pc_plus_4_D~13_combout ;
wire \pc_plus_4_D~14_combout ;
wire \pc_plus_4_D~15_combout ;
wire \pc_plus_4_D~17_combout ;
wire \pc_plus_4_D~19_combout ;
wire \pc_plus_4_D~20_combout ;
wire \pc_plus_4_D~23_combout ;
wire \pc_plus_4_D~25_combout ;
wire \pc_plus_4_D~27_combout ;
wire \pc_plus_4_D~28_combout ;
wire \pc_plus_4_D~29_combout ;
wire \pc_plus_4_D~30_combout ;
wire \portB~112_combout ;
wire \portB~113_combout ;
wire \portB~114_combout ;
wire \portB~116_combout ;
wire \portA~70_combout ;
wire \portA~71_combout ;
wire \portA~72_combout ;
wire \comb~3_combout ;
wire \PROGRAM_COUNTER|pc_out[10]~31_combout ;
wire \ALU|ShiftRight0~91_combout ;
wire \btbframes.frameblocks[2].tag[27]~3_combout ;
wire \btbframes.frameblocks[0].tag[27]~3_combout ;
wire \always3~3_combout ;
wire \btbframes.frameblocks[2].valid~2_combout ;
wire \btbframes.frameblocks[1].valid~2_combout ;
wire \btbframes.frameblocks[3].valid~2_combout ;
wire \jal_EX~2_combout ;
wire \instruction_D~70_combout ;
wire \instruction_D~71_combout ;
wire \instruction_D~72_combout ;
wire \instruction_D~73_combout ;
wire \instruction_D~75_combout ;
wire \instruction_D~77_combout ;
wire \instruction_D~78_combout ;
wire \instruction_D~79_combout ;
wire \instruction_D~92_combout ;
wire \btbframes.frameblocks[1].jump_add[3]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[3]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[4]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[6]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[7]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[8]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[10]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[10]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[11]~feeder_combout ;
wire \btbframes.frameblocks[0].jump_add[11]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[12]~feeder_combout ;
wire \btbframes.frameblocks[0].jump_add[13]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[13]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[14]~feeder_combout ;
wire \btbframes.frameblocks[0].jump_add[14]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[15]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[16]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[16]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[18]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[19]~feeder_combout ;
wire \btbframes.frameblocks[0].jump_add[20]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[21]~feeder_combout ;
wire \btbframes.frameblocks[3].jump_add[21]~feeder_combout ;
wire \btbframes.frameblocks[3].jump_add[23]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[23]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[24]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[26]~feeder_combout ;
wire \btbframes.frameblocks[3].jump_add[26]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[28]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[28]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[30]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[31]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[0]~feeder_combout ;
wire \btbframes.frameblocks[0].tag[1]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[2]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[3]~feeder_combout ;
wire \btbframes.frameblocks[0].tag[3]~feeder_combout ;
wire \btbframes.frameblocks[2].tag[5]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[8]~feeder_combout ;
wire \btbframes.frameblocks[1].tag[9]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[9]~feeder_combout ;
wire \btbframes.frameblocks[1].tag[15]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[15]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[16]~feeder_combout ;
wire \btbframes.frameblocks[2].tag[16]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[18]~feeder_combout ;
wire \btbframes.frameblocks[1].tag[18]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[20]~feeder_combout ;
wire \btbframes.frameblocks[2].tag[20]~feeder_combout ;
wire \btbframes.frameblocks[0].tag[21]~feeder_combout ;
wire \btbframes.frameblocks[2].tag[22]~feeder_combout ;
wire \btbframes.frameblocks[1].tag[23]~feeder_combout ;
wire \btbframes.frameblocks[0].tag[24]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[26]~feeder_combout ;
wire \btbframes.frameblocks[2].tag[26]~feeder_combout ;
wire \btbframes.frameblocks[3].tag[27]~feeder_combout ;
wire \dmemload_WB[4]~feeder_combout ;
wire \dmemload_WB[15]~feeder_combout ;
wire \dmemload_WB[18]~feeder_combout ;
wire \dmemload_WB[19]~feeder_combout ;
wire \btbframes.frameblocks[2].jump_add[1]~feeder_combout ;
wire \btbframes.frameblocks[1].jump_add[0]~feeder_combout ;
wire \pc_plus_4_WB[18]~feeder_combout ;
wire \instruction_D~68_combout ;
wire \ALUSrc_EX~0_combout ;
wire \instruction_D~69_combout ;
wire \instruction_D~66_combout ;
wire \instruction_D~67_combout ;
wire \j_EX~3_combout ;
wire \j_EX~2_combout ;
wire \j_EX~q ;
wire \predicted_M~3_combout ;
wire \j_M~0_combout ;
wire \j_M~q ;
wire \en_EX~0_combout ;
wire \wsel_M~0_combout ;
wire \jal_M~0_combout ;
wire \jal_M~q ;
wire \branch_or_jump~0_combout ;
wire \predicted_M~2_combout ;
wire \predicted_M~q ;
wire \beq_M~0_combout ;
wire \always4~3_combout ;
wire \beq_M~q ;
wire \zero_M~7_combout ;
wire \zero_M~8_combout ;
wire \zero_M~9_combout ;
wire \zero_M~10_combout ;
wire \zero_M~11_combout ;
wire \zero_M~0_combout ;
wire \zero_M~1_combout ;
wire \zero_M~2_combout ;
wire \zero_M~3_combout ;
wire \zero_M~4_combout ;
wire \zero_M~6_combout ;
wire \zero_M~12_combout ;
wire \zero_M~q ;
wire \branch_taken~0_combout ;
wire \branch_or_jump~1_combout ;
wire \pc_plus_4_D~1_combout ;
wire \branch_or_jump~2_combout ;
wire \pc_plus_4_EX~1_combout ;
wire \pc_plus_4_M~1_combout ;
wire \pc_plus_4_WB[0]~feeder_combout ;
wire \halt_M~0_combout ;
wire \halt_M~q ;
wire \halt_WB~_Duplicate_1_q ;
wire \always4~2_combout ;
wire \lui_M~0_combout ;
wire \lui_M~q ;
wire \lui_WB~q ;
wire \jal_WB~feeder_combout ;
wire \jal_WB~q ;
wire \wdat_WB[0]~60_combout ;
wire \wdat_WB[0]~61_combout ;
wire \instruction_D~65_combout ;
wire \instruction_D~64_combout ;
wire \dWEN_EX~0_combout ;
wire \dWEN_EX~q ;
wire \rdata2_M[16]~0_combout ;
wire \rdata2_M[16]~1_combout ;
wire \sw_forwarding_output~27_combout ;
wire \rdata2_M~2_combout ;
wire \rdata2_M~3_combout ;
wire \sw_forwarding_output~28_combout ;
wire \lui_EX~0_combout ;
wire \MemToReg_EX~2_combout ;
wire \MemToReg_EX~q ;
wire \memToReg_M~0_combout ;
wire \memToReg_M~q ;
wire \memToReg_WB~q ;
wire \wdat_WB[1]~58_combout ;
wire \pc_plus_4_M~0_combout ;
wire \wdat_WB[1]~59_combout ;
wire \rdata2_M~4_combout ;
wire \rdata2_M~5_combout ;
wire \pc_plus_4[2]~0_combout ;
wire \pc_plus_4_D~3_combout ;
wire \pc_plus_4_EX~3_combout ;
wire \pc_plus_4_M~3_combout ;
wire \wdat_WB[2]~56_combout ;
wire \wdat_WB[2]~57_combout ;
wire \Equal2~0_combout ;
wire \instruction_D~91_combout ;
wire \imm_EX~5_combout ;
wire \instruction_D~83_combout ;
wire \instruction_D~80_combout ;
wire \instruction_D~82_combout ;
wire \ShiftOp_EX~0_combout ;
wire \instruction_D~85_combout ;
wire \ShiftOp_EX~1_combout ;
wire \ShiftOp_EX~q ;
wire \portB~88_combout ;
wire \portB~93_combout ;
wire \portB~98_combout ;
wire \portB~99_combout ;
wire \portB~100_combout ;
wire \rdata2_EX~58_combout ;
wire \rdata2_EX~59_combout ;
wire \Equal3~2_combout ;
wire \rdata1_EX[15]~0_combout ;
wire \always2~2_combout ;
wire \rdata1_EX[15]~1_combout ;
wire \rdata2_M~6_combout ;
wire \rdata2_M~7_combout ;
wire \pc_plus_4_EX~2_combout ;
wire \pc_plus_4_M~2_combout ;
wire \wdat_WB[3]~64_combout ;
wire \wdat_WB[3]~65_combout ;
wire \rdata2_M~8_combout ;
wire \sw_forwarding_output~30_combout ;
wire \rdata2_M~9_combout ;
wire \portB~104_combout ;
wire \imm_EX~15_combout ;
wire \portB~105_combout ;
wire \instruction_D~93_combout ;
wire \imm_EX~7_combout ;
wire \portB~106_combout ;
wire \portB~107_combout ;
wire \instruction_D~74_combout ;
wire \rdata2_EX~62_combout ;
wire \rdata2_EX~63_combout ;
wire \rdata2_M~10_combout ;
wire \pc_plus_4_EX~5_combout ;
wire \pc_plus_4_M~5_combout ;
wire \wdat_WB[4]~63_combout ;
wire \rdata2_M~11_combout ;
wire \pc_plus_4_EX~4_combout ;
wire \pc_plus_4_M~4_combout ;
wire \wdat_WB[5]~54_combout ;
wire \wdat_WB[5]~55_combout ;
wire \sw_forwarding_output~26_combout ;
wire \rdata2_M~12_combout ;
wire \rdata2_M~13_combout ;
wire \pc_plus_4_EX~7_combout ;
wire \pc_plus_4_M~7_combout ;
wire \wdat_WB[6]~52_combout ;
wire \wdat_WB[6]~53_combout ;
wire \instruction_D~95_combout ;
wire \imm_EX~9_combout ;
wire \portB~14_combout ;
wire \portB~83_combout ;
wire \portB~115_combout ;
wire \portB~84_combout ;
wire \rdata2_EX~50_combout ;
wire \rdata2_EX~51_combout ;
wire \rdata2_M~14_combout ;
wire \rdata2_M~15_combout ;
wire \sw_forwarding_output~24_combout ;
wire \pc_plus_4[2]~1 ;
wire \pc_plus_4[3]~3 ;
wire \pc_plus_4[4]~5 ;
wire \pc_plus_4[5]~7 ;
wire \pc_plus_4[6]~9 ;
wire \pc_plus_4[7]~10_combout ;
wire \pc_plus_4_D~6_combout ;
wire \pc_plus_4_EX~6_combout ;
wire \pc_plus_4_M~6_combout ;
wire \dmemload_WB[7]~feeder_combout ;
wire \wdat_WB[7]~50_combout ;
wire \wdat_WB[7]~51_combout ;
wire \rdata2_M~16_combout ;
wire \rdata2_M~17_combout ;
wire \pc_plus_4_M~9_combout ;
wire \wdat_WB[8]~44_combout ;
wire \wdat_WB[8]~45_combout ;
wire \sw_forwarding_output~21_combout ;
wire \rdata2_M~18_combout ;
wire \rdata2_M~19_combout ;
wire \pc_plus_4_EX~8_combout ;
wire \pc_plus_4_M~8_combout ;
wire \dmemload_WB[9]~feeder_combout ;
wire \wdat_WB[9]~42_combout ;
wire \wdat_WB[9]~43_combout ;
wire \sw_forwarding_output~20_combout ;
wire \instruction_D~90_combout ;
wire \imm_EX~4_combout ;
wire \portB~71_combout ;
wire \portB~72_combout ;
wire \portB~73_combout ;
wire \rdata2_EX~40_combout ;
wire \rdata2_EX~41_combout ;
wire \rdata2_M~20_combout ;
wire \rdata2_M~21_combout ;
wire \pc_plus_4_EX~11_combout ;
wire \pc_plus_4_M~11_combout ;
wire \wdat_WB[10]~48_combout ;
wire \wdat_WB[10]~49_combout ;
wire \sw_forwarding_output~23_combout ;
wire \rdata2_M~22_combout ;
wire \rdata2_M~23_combout ;
wire \sw_forwarding_output~22_combout ;
wire \pc_plus_4_EX~10_combout ;
wire \pc_plus_4_M~10_combout ;
wire \wdat_WB[11]~46_combout ;
wire \wdat_WB[11]~47_combout ;
wire \rdata2_M~24_combout ;
wire \rdata2_M~25_combout ;
wire \rdata2_EX~38_combout ;
wire \rdata2_EX~39_combout ;
wire \sw_forwarding_output~19_combout ;
wire \rdata2_M~26_combout ;
wire \wdat_WB[12]~40_combout ;
wire \pc_plus_4_M~13_combout ;
wire \wdat_WB[12]~41_combout ;
wire \rdata2_M~27_combout ;
wire \sw_forwarding_output~18_combout ;
wire \pc_plus_4_EX~12_combout ;
wire \pc_plus_4_M~12_combout ;
wire \wdat_WB[13]~38_combout ;
wire \wdat_WB[13]~39_combout ;
wire \rdata2_M~28_combout ;
wire \rdata2_M~29_combout ;
wire \instruction_D~87_combout ;
wire \imm_EX~1_combout ;
wire \portB~65_combout ;
wire \portB~111_combout ;
wire \portB~66_combout ;
wire \rdata2_EX~34_combout ;
wire \rdata2_EX~35_combout ;
wire \rdata2_M~30_combout ;
wire \pc_plus_4_M~15_combout ;
wire \wdat_WB[14]~36_combout ;
wire \wdat_WB[14]~37_combout ;
wire \rdata2_M~31_combout ;
wire \pc_plus_4_M~14_combout ;
wire \wdat_WB[15]~34_combout ;
wire \wdat_WB[15]~35_combout ;
wire \instruction_D~86_combout ;
wire \imm_EX~0_combout ;
wire \portB~63_combout ;
wire \portB~110_combout ;
wire \portB~64_combout ;
wire \rdata2_EX~32_combout ;
wire \rdata2_EX~33_combout ;
wire \rdata2_M~32_combout ;
wire \sw_forwarding_output~16_combout ;
wire \rdata2_M~33_combout ;
wire \instruction_D~81_combout ;
wire \imm_EX~11_combout ;
wire \imm_M~15_combout ;
wire \wdat_WB[28]~1_combout ;
wire \wdat_WB[28]~0_combout ;
wire \wdat_WB[16]~32_combout ;
wire \wdat_WB[16]~33_combout ;
wire \sw_forwarding_output~15_combout ;
wire \rdata2_EX~30_combout ;
wire \portB~61_combout ;
wire \portB~62_combout ;
wire \rdata2_EX~31_combout ;
wire \rdata2_M~34_combout ;
wire \rdata2_M~35_combout ;
wire \pc_plus_4[7]~11 ;
wire \pc_plus_4[8]~13 ;
wire \pc_plus_4[9]~15 ;
wire \pc_plus_4[10]~17 ;
wire \pc_plus_4[11]~19 ;
wire \pc_plus_4[12]~21 ;
wire \pc_plus_4[13]~23 ;
wire \pc_plus_4[14]~25 ;
wire \pc_plus_4[15]~27 ;
wire \pc_plus_4[16]~29 ;
wire \pc_plus_4[17]~30_combout ;
wire \pc_plus_4_D~16_combout ;
wire \pc_plus_4_EX~16_combout ;
wire \pc_plus_4_M~16_combout ;
wire \wdat_WB[17]~30_combout ;
wire \wdat_WB[17]~31_combout ;
wire \instruction_D~84_combout ;
wire \imm_EX~12_combout ;
wire \imm_M~14_combout ;
wire \sw_forwarding_output~14_combout ;
wire \rdata2_EX~28_combout ;
wire \rdata2_EX~29_combout ;
wire \rdata2_M~36_combout ;
wire \rdata2_M~37_combout ;
wire \imm_EX~13_combout ;
wire \imm_M~13_combout ;
wire \wdat_WB[18]~28_combout ;
wire \wdat_WB[18]~29_combout ;
wire \sw_forwarding_output~13_combout ;
wire \portB~55_combout ;
wire \portB~54_combout ;
wire \portB~56_combout ;
wire \rdata2_EX~26_combout ;
wire \rdata2_EX~27_combout ;
wire \rdata2_M~38_combout ;
wire \rdata2_M~39_combout ;
wire \imm_EX~14_combout ;
wire \imm_M~12_combout ;
wire \sw_forwarding_output~12_combout ;
wire \imm_WB[3]~feeder_combout ;
wire \pc_plus_4[17]~31 ;
wire \pc_plus_4[18]~33 ;
wire \pc_plus_4[19]~34_combout ;
wire \pc_plus_4_D~18_combout ;
wire \pc_plus_4_EX~18_combout ;
wire \pc_plus_4_M~18_combout ;
wire \wdat_WB[19]~26_combout ;
wire \wdat_WB[19]~27_combout ;
wire \portB~51_combout ;
wire \portB~52_combout ;
wire \portB~53_combout ;
wire \rdata2_EX~24_combout ;
wire \rdata2_EX~25_combout ;
wire \rdata2_M~40_combout ;
wire \rdata2_M~41_combout ;
wire \sw_forwarding_output~11_combout ;
wire \rdata2_M~42_combout ;
wire \imm_M~11_combout ;
wire \pc_plus_4[19]~35 ;
wire \pc_plus_4[20]~36_combout ;
wire \pc_plus_4_D~21_combout ;
wire \pc_plus_4_EX~21_combout ;
wire \pc_plus_4_M~21_combout ;
wire \pc_plus_4_WB[20]~feeder_combout ;
wire \wdat_WB[20]~24_combout ;
wire \wdat_WB[20]~25_combout ;
wire \rdata2_M~43_combout ;
wire \sw_forwarding_output~10_combout ;
wire \imm_EX~10_combout ;
wire \imm_M~10_combout ;
wire \wdat_WB[21]~22_combout ;
wire \wdat_WB[21]~23_combout ;
wire \ExtOp_EX~1_combout ;
wire \ExtOp_EX~q ;
wire \sign_ext[16]~0_combout ;
wire \portB~45_combout ;
wire \portB~46_combout ;
wire \portB~47_combout ;
wire \rdata2_EX~20_combout ;
wire \rdata2_EX~21_combout ;
wire \rdata2_M~44_combout ;
wire \rdata2_M~45_combout ;
wire \rdata2_EX~18_combout ;
wire \rdata2_EX~19_combout ;
wire \rdata2_M~46_combout ;
wire \imm_M~9_combout ;
wire \imm_WB[6]~feeder_combout ;
wire \pc_plus_4_M~23_combout ;
wire \pc_plus_4_WB[22]~feeder_combout ;
wire \wdat_WB[22]~20_combout ;
wire \wdat_WB[22]~21_combout ;
wire \rdata2_M~47_combout ;
wire \instruction_D~94_combout ;
wire \imm_EX~8_combout ;
wire \imm_M~8_combout ;
wire \sw_forwarding_output~8_combout ;
wire \pc_plus_4[20]~37 ;
wire \pc_plus_4[21]~39 ;
wire \pc_plus_4[22]~41 ;
wire \pc_plus_4[23]~42_combout ;
wire \pc_plus_4_D~22_combout ;
wire \pc_plus_4_EX~22_combout ;
wire \pc_plus_4_M~22_combout ;
wire \wdat_WB[23]~18_combout ;
wire \wdat_WB[23]~19_combout ;
wire \rdata2_EX~16_combout ;
wire \rdata2_EX~17_combout ;
wire \rdata2_M~48_combout ;
wire \rdata2_M~49_combout ;
wire \imm_M~7_combout ;
wire \pc_plus_4_EX~25_combout ;
wire \pc_plus_4_M~25_combout ;
wire \wdat_WB[24]~16_combout ;
wire \wdat_WB[24]~17_combout ;
wire \rdata2_EX~14_combout ;
wire \rdata2_EX~15_combout ;
wire \sw_forwarding_output~7_combout ;
wire \rdata2_M~50_combout ;
wire \rdata2_M~51_combout ;
wire \imm_M~6_combout ;
wire \imm_WB[9]~feeder_combout ;
wire \pc_plus_4[23]~43 ;
wire \pc_plus_4[24]~45 ;
wire \pc_plus_4[25]~46_combout ;
wire \pc_plus_4_D~24_combout ;
wire \pc_plus_4_EX~24_combout ;
wire \pc_plus_4_M~24_combout ;
wire \wdat_WB[25]~14_combout ;
wire \wdat_WB[25]~15_combout ;
wire \sw_forwarding_output~6_combout ;
wire \rdata2_M~52_combout ;
wire \rdata2_M~53_combout ;
wire \imm_M~5_combout ;
wire \pc_plus_4_EX~27_combout ;
wire \pc_plus_4_M~27_combout ;
wire \wdat_WB[26]~12_combout ;
wire \wdat_WB[26]~13_combout ;
wire \portB~30_combout ;
wire \portB~31_combout ;
wire \portB~32_combout ;
wire \rdata2_EX~10_combout ;
wire \rdata2_EX~11_combout ;
wire \rdata2_M~54_combout ;
wire \rdata2_M~55_combout ;
wire \pc_plus_4[25]~47 ;
wire \pc_plus_4[26]~49 ;
wire \pc_plus_4[27]~50_combout ;
wire \pc_plus_4_D~26_combout ;
wire \pc_plus_4_EX~26_combout ;
wire \pc_plus_4_M~26_combout ;
wire \wdat_WB[27]~10_combout ;
wire \wdat_WB[27]~11_combout ;
wire \imm_M~4_combout ;
wire \sw_forwarding_output~4_combout ;
wire \rdata2_M~56_combout ;
wire \rdata2_M~57_combout ;
wire \wdat_WB[28]~8_combout ;
wire \instruction_D~89_combout ;
wire \imm_EX~3_combout ;
wire \imm_M~3_combout ;
wire \wdat_WB[28]~9_combout ;
wire \portB~24_combout ;
wire \portB~25_combout ;
wire \portB~26_combout ;
wire \rdata2_EX~6_combout ;
wire \rdata2_EX~7_combout ;
wire \sw_forwarding_output~3_combout ;
wire \rdata2_M~58_combout ;
wire \rdata2_M~59_combout ;
wire \instruction_D~88_combout ;
wire \imm_EX~2_combout ;
wire \imm_M~2_combout ;
wire \sw_forwarding_output~2_combout ;
wire \imm_WB[13]~feeder_combout ;
wire \pc_plus_4_M~28_combout ;
wire \wdat_WB[29]~6_combout ;
wire \wdat_WB[29]~7_combout ;
wire \portB~21_combout ;
wire \portB~22_combout ;
wire \portB~23_combout ;
wire \rdata2_EX~4_combout ;
wire \rdata2_EX~5_combout ;
wire \rdata2_M~60_combout ;
wire \rdata2_M~61_combout ;
wire \imm_M~1_combout ;
wire \pc_plus_4[27]~51 ;
wire \pc_plus_4[28]~53 ;
wire \pc_plus_4[29]~55 ;
wire \pc_plus_4[30]~56_combout ;
wire \pc_plus_4_D~31_combout ;
wire \pc_plus_4_EX~31_combout ;
wire \pc_plus_4_M~31_combout ;
wire \pc_plus_4_WB[30]~feeder_combout ;
wire \wdat_WB[30]~4_combout ;
wire \wdat_WB[30]~5_combout ;
wire \sw_forwarding_output~1_combout ;
wire \portB~18_combout ;
wire \portB~19_combout ;
wire \portB~20_combout ;
wire \rdata2_EX~2_combout ;
wire \rdata2_EX~3_combout ;
wire \rdata2_M~62_combout ;
wire \rdata2_M~63_combout ;
wire \imm_M~0_combout ;
wire \imm_WB[15]~feeder_combout ;
wire \pc_plus_4_EX~30_combout ;
wire \pc_plus_4_M~30_combout ;
wire \wdat_WB[31]~2_combout ;
wire \wdat_WB[31]~3_combout ;
wire \sw_forwarding_output~0_combout ;
wire \rdata2_EX~0_combout ;
wire \rdata2_EX~1_combout ;
wire \rdata2_M~64_combout ;
wire \rdata2_M~65_combout ;
wire \porto_M~4_combout ;
wire \dWEN_M~0_combout ;
wire \dREN_EX~0_combout ;
wire \dREN_EX~1_combout ;
wire \dREN_EX~q ;
wire \dREN_M~0_combout ;
wire \instruction_D~76_combout ;
wire \instruction_EX~6_combout ;
wire \rdata1_EX~64_combout ;
wire \rdata1_EX~65_combout ;
wire \regWrite_M~0_combout ;
wire \regWrite_M~q ;
wire \regWrite_WB~q ;
wire \portA~68_combout ;
wire \portA~73_combout ;
wire \portA~69_combout ;
wire \porto_M~35_combout ;
wire \porto_M~5_combout ;
wire \porto_M~6_combout ;
wire \porto_M~7_combout ;
wire \porto_M~8_combout ;
wire \porto_M~36_combout ;
wire \porto_M~9_combout ;
wire \porto_M~10_combout ;
wire \porto_M~11_combout ;
wire \porto_M~12_combout ;
wire \porto_M~13_combout ;
wire \porto_M~14_combout ;
wire \porto_M~15_combout ;
wire \porto_M~16_combout ;
wire \porto_M~17_combout ;
wire \porto_M~18_combout ;
wire \porto_M~19_combout ;
wire \porto_M~20_combout ;
wire \porto_M~21_combout ;
wire \porto_M~22_combout ;
wire \porto_M~23_combout ;
wire \porto_M~24_combout ;
wire \porto_M~25_combout ;
wire \porto_M~26_combout ;
wire \porto_M~27_combout ;
wire \porto_M~28_combout ;
wire \porto_M~29_combout ;
wire \porto_M~30_combout ;
wire \porto_M~31_combout ;
wire \porto_M~32_combout ;
wire \porto_M~33_combout ;
wire \porto_M~34_combout ;
wire [4:0] wsel_WB;
wire [4:0] wsel_M;
wire [31:0] rdata2_EX;
wire [31:0] rdata1_M;
wire [31:0] rdata1_EX;
wire [31:0] porto_WB;
wire [31:0] pc_plus_4_WB;
wire [31:0] pc_plus_4_M;
wire [31:0] pc_plus_4_EX;
wire [31:0] pc_plus_4_D;
wire [5:0] op_EX;
wire [5:0] op_D;
wire [31:0] instruction_M;
wire [31:0] instruction_EX;
wire [31:0] instruction_D;
wire [15:0] imm_WB;
wire [15:0] imm_M;
wire [15:0] imm_EX;
wire [31:0] dmemload_WB;
wire [27:0] \btbframes.frameblocks[3].tag ;
wire [31:0] \btbframes.frameblocks[3].jump_add ;
wire [1:0] \btbframes.frameblocks[3].curr_state ;
wire [27:0] \btbframes.frameblocks[2].tag ;
wire [31:0] \btbframes.frameblocks[2].jump_add ;
wire [1:0] \btbframes.frameblocks[2].curr_state ;
wire [27:0] \btbframes.frameblocks[1].tag ;
wire [31:0] \btbframes.frameblocks[1].jump_add ;
wire [1:0] \btbframes.frameblocks[1].curr_state ;
wire [27:0] \btbframes.frameblocks[0].tag ;
wire [31:0] \btbframes.frameblocks[0].jump_add ;
wire [1:0] \btbframes.frameblocks[0].curr_state ;
wire [3:0] ALUOp_EX;


btb BTB(
	.pc_out_3(pc_out_3),
	.pc_out_2(pc_out_2),
	.pc_out_5(pc_out_5),
	.pc_out_4(pc_out_4),
	.pc_out_7(pc_out_7),
	.pc_out_6(pc_out_6),
	.pc_out_9(pc_out_9),
	.pc_out_8(pc_out_8),
	.pc_out_11(pc_out_11),
	.pc_out_10(pc_out_10),
	.pc_out_13(pc_out_13),
	.pc_out_12(pc_out_12),
	.pc_out_15(pc_out_15),
	.pc_out_14(pc_out_14),
	.pc_out_17(pc_out_17),
	.pc_out_16(pc_out_16),
	.pc_out_19(pc_out_19),
	.pc_out_18(pc_out_18),
	.pc_out_21(pc_out_21),
	.pc_out_20(pc_out_20),
	.pc_out_23(pc_out_23),
	.pc_out_22(pc_out_22),
	.pc_out_25(pc_out_25),
	.pc_out_24(pc_out_24),
	.pc_out_27(pc_out_27),
	.pc_out_26(pc_out_26),
	.pc_out_29(pc_out_29),
	.pc_out_28(pc_out_28),
	.pc_out_31(pc_out_31),
	.pc_out_30(pc_out_30),
	.btbframesframeblocks2tag_1(\btbframes.frameblocks[2].tag [1]),
	.btbframesframeblocks1tag_1(\btbframes.frameblocks[1].tag [1]),
	.btbframesframeblocks0tag_1(\btbframes.frameblocks[0].tag [1]),
	.btbframesframeblocks3tag_1(\btbframes.frameblocks[3].tag [1]),
	.btbframesframeblocks1tag_0(\btbframes.frameblocks[1].tag [0]),
	.btbframesframeblocks2tag_0(\btbframes.frameblocks[2].tag [0]),
	.btbframesframeblocks0tag_0(\btbframes.frameblocks[0].tag [0]),
	.btbframesframeblocks3tag_0(\btbframes.frameblocks[3].tag [0]),
	.btbframesframeblocks2tag_3(\btbframes.frameblocks[2].tag [3]),
	.btbframesframeblocks1tag_3(\btbframes.frameblocks[1].tag [3]),
	.btbframesframeblocks0tag_3(\btbframes.frameblocks[0].tag [3]),
	.btbframesframeblocks3tag_3(\btbframes.frameblocks[3].tag [3]),
	.btbframesframeblocks1tag_2(\btbframes.frameblocks[1].tag [2]),
	.btbframesframeblocks2tag_2(\btbframes.frameblocks[2].tag [2]),
	.btbframesframeblocks0tag_2(\btbframes.frameblocks[0].tag [2]),
	.btbframesframeblocks3tag_2(\btbframes.frameblocks[3].tag [2]),
	.btbframesframeblocks2tag_5(\btbframes.frameblocks[2].tag [5]),
	.btbframesframeblocks1tag_5(\btbframes.frameblocks[1].tag [5]),
	.btbframesframeblocks0tag_5(\btbframes.frameblocks[0].tag [5]),
	.btbframesframeblocks3tag_5(\btbframes.frameblocks[3].tag [5]),
	.btbframesframeblocks1tag_4(\btbframes.frameblocks[1].tag [4]),
	.btbframesframeblocks2tag_4(\btbframes.frameblocks[2].tag [4]),
	.btbframesframeblocks0tag_4(\btbframes.frameblocks[0].tag [4]),
	.btbframesframeblocks3tag_4(\btbframes.frameblocks[3].tag [4]),
	.btbframesframeblocks2tag_7(\btbframes.frameblocks[2].tag [7]),
	.btbframesframeblocks1tag_7(\btbframes.frameblocks[1].tag [7]),
	.btbframesframeblocks0tag_7(\btbframes.frameblocks[0].tag [7]),
	.btbframesframeblocks3tag_7(\btbframes.frameblocks[3].tag [7]),
	.btbframesframeblocks1tag_6(\btbframes.frameblocks[1].tag [6]),
	.btbframesframeblocks2tag_6(\btbframes.frameblocks[2].tag [6]),
	.btbframesframeblocks0tag_6(\btbframes.frameblocks[0].tag [6]),
	.btbframesframeblocks3tag_6(\btbframes.frameblocks[3].tag [6]),
	.btbframesframeblocks2tag_9(\btbframes.frameblocks[2].tag [9]),
	.btbframesframeblocks1tag_9(\btbframes.frameblocks[1].tag [9]),
	.btbframesframeblocks0tag_9(\btbframes.frameblocks[0].tag [9]),
	.btbframesframeblocks3tag_9(\btbframes.frameblocks[3].tag [9]),
	.btbframesframeblocks1tag_8(\btbframes.frameblocks[1].tag [8]),
	.btbframesframeblocks2tag_8(\btbframes.frameblocks[2].tag [8]),
	.btbframesframeblocks0tag_8(\btbframes.frameblocks[0].tag [8]),
	.btbframesframeblocks3tag_8(\btbframes.frameblocks[3].tag [8]),
	.btbframesframeblocks2tag_11(\btbframes.frameblocks[2].tag [11]),
	.btbframesframeblocks1tag_11(\btbframes.frameblocks[1].tag [11]),
	.btbframesframeblocks0tag_11(\btbframes.frameblocks[0].tag [11]),
	.btbframesframeblocks3tag_11(\btbframes.frameblocks[3].tag [11]),
	.btbframesframeblocks1tag_10(\btbframes.frameblocks[1].tag [10]),
	.btbframesframeblocks2tag_10(\btbframes.frameblocks[2].tag [10]),
	.btbframesframeblocks0tag_10(\btbframes.frameblocks[0].tag [10]),
	.btbframesframeblocks3tag_10(\btbframes.frameblocks[3].tag [10]),
	.btbframesframeblocks2tag_13(\btbframes.frameblocks[2].tag [13]),
	.btbframesframeblocks1tag_13(\btbframes.frameblocks[1].tag [13]),
	.btbframesframeblocks0tag_13(\btbframes.frameblocks[0].tag [13]),
	.btbframesframeblocks3tag_13(\btbframes.frameblocks[3].tag [13]),
	.btbframesframeblocks1tag_12(\btbframes.frameblocks[1].tag [12]),
	.btbframesframeblocks2tag_12(\btbframes.frameblocks[2].tag [12]),
	.btbframesframeblocks0tag_12(\btbframes.frameblocks[0].tag [12]),
	.btbframesframeblocks3tag_12(\btbframes.frameblocks[3].tag [12]),
	.btbframesframeblocks2tag_15(\btbframes.frameblocks[2].tag [15]),
	.btbframesframeblocks1tag_15(\btbframes.frameblocks[1].tag [15]),
	.btbframesframeblocks0tag_15(\btbframes.frameblocks[0].tag [15]),
	.btbframesframeblocks3tag_15(\btbframes.frameblocks[3].tag [15]),
	.btbframesframeblocks1tag_14(\btbframes.frameblocks[1].tag [14]),
	.btbframesframeblocks2tag_14(\btbframes.frameblocks[2].tag [14]),
	.btbframesframeblocks0tag_14(\btbframes.frameblocks[0].tag [14]),
	.btbframesframeblocks3tag_14(\btbframes.frameblocks[3].tag [14]),
	.btbframesframeblocks2tag_17(\btbframes.frameblocks[2].tag [17]),
	.btbframesframeblocks1tag_17(\btbframes.frameblocks[1].tag [17]),
	.btbframesframeblocks0tag_17(\btbframes.frameblocks[0].tag [17]),
	.btbframesframeblocks3tag_17(\btbframes.frameblocks[3].tag [17]),
	.btbframesframeblocks1tag_16(\btbframes.frameblocks[1].tag [16]),
	.btbframesframeblocks2tag_16(\btbframes.frameblocks[2].tag [16]),
	.btbframesframeblocks0tag_16(\btbframes.frameblocks[0].tag [16]),
	.btbframesframeblocks3tag_16(\btbframes.frameblocks[3].tag [16]),
	.btbframesframeblocks2tag_19(\btbframes.frameblocks[2].tag [19]),
	.btbframesframeblocks1tag_19(\btbframes.frameblocks[1].tag [19]),
	.btbframesframeblocks0tag_19(\btbframes.frameblocks[0].tag [19]),
	.btbframesframeblocks3tag_19(\btbframes.frameblocks[3].tag [19]),
	.btbframesframeblocks1tag_18(\btbframes.frameblocks[1].tag [18]),
	.btbframesframeblocks2tag_18(\btbframes.frameblocks[2].tag [18]),
	.btbframesframeblocks0tag_18(\btbframes.frameblocks[0].tag [18]),
	.btbframesframeblocks3tag_18(\btbframes.frameblocks[3].tag [18]),
	.btbframesframeblocks2tag_21(\btbframes.frameblocks[2].tag [21]),
	.btbframesframeblocks1tag_21(\btbframes.frameblocks[1].tag [21]),
	.btbframesframeblocks0tag_21(\btbframes.frameblocks[0].tag [21]),
	.btbframesframeblocks3tag_21(\btbframes.frameblocks[3].tag [21]),
	.btbframesframeblocks1tag_20(\btbframes.frameblocks[1].tag [20]),
	.btbframesframeblocks2tag_20(\btbframes.frameblocks[2].tag [20]),
	.btbframesframeblocks0tag_20(\btbframes.frameblocks[0].tag [20]),
	.btbframesframeblocks3tag_20(\btbframes.frameblocks[3].tag [20]),
	.btbframesframeblocks2tag_23(\btbframes.frameblocks[2].tag [23]),
	.btbframesframeblocks1tag_23(\btbframes.frameblocks[1].tag [23]),
	.btbframesframeblocks0tag_23(\btbframes.frameblocks[0].tag [23]),
	.btbframesframeblocks3tag_23(\btbframes.frameblocks[3].tag [23]),
	.btbframesframeblocks1tag_22(\btbframes.frameblocks[1].tag [22]),
	.btbframesframeblocks2tag_22(\btbframes.frameblocks[2].tag [22]),
	.btbframesframeblocks0tag_22(\btbframes.frameblocks[0].tag [22]),
	.btbframesframeblocks3tag_22(\btbframes.frameblocks[3].tag [22]),
	.btbframesframeblocks2tag_25(\btbframes.frameblocks[2].tag [25]),
	.btbframesframeblocks1tag_25(\btbframes.frameblocks[1].tag [25]),
	.btbframesframeblocks0tag_25(\btbframes.frameblocks[0].tag [25]),
	.btbframesframeblocks3tag_25(\btbframes.frameblocks[3].tag [25]),
	.btbframesframeblocks1tag_24(\btbframes.frameblocks[1].tag [24]),
	.btbframesframeblocks2tag_24(\btbframes.frameblocks[2].tag [24]),
	.btbframesframeblocks0tag_24(\btbframes.frameblocks[0].tag [24]),
	.btbframesframeblocks3tag_24(\btbframes.frameblocks[3].tag [24]),
	.btbframesframeblocks2tag_27(\btbframes.frameblocks[2].tag [27]),
	.btbframesframeblocks1tag_27(\btbframes.frameblocks[1].tag [27]),
	.btbframesframeblocks0tag_27(\btbframes.frameblocks[0].tag [27]),
	.btbframesframeblocks3tag_27(\btbframes.frameblocks[3].tag [27]),
	.btbframesframeblocks1tag_26(\btbframes.frameblocks[1].tag [26]),
	.btbframesframeblocks2tag_26(\btbframes.frameblocks[2].tag [26]),
	.btbframesframeblocks0tag_26(\btbframes.frameblocks[0].tag [26]),
	.btbframesframeblocks3tag_26(\btbframes.frameblocks[3].tag [26]),
	.btbframesframeblocks2valid(\btbframes.frameblocks[2].valid~q ),
	.btbframesframeblocks1valid(\btbframes.frameblocks[1].valid~q ),
	.btbframesframeblocks0valid(\btbframes.frameblocks[0].valid~q ),
	.btbframesframeblocks3valid(\btbframes.frameblocks[3].valid~q ),
	.btbframesframeblocks1curr_state_1(\btbframes.frameblocks[1].curr_state [1]),
	.btbframesframeblocks2curr_state_1(\btbframes.frameblocks[2].curr_state [1]),
	.btbframesframeblocks0curr_state_1(\btbframes.frameblocks[0].curr_state [1]),
	.btbframesframeblocks3curr_state_1(\btbframes.frameblocks[3].curr_state [1]),
	.predicted(\BTB|predicted~18_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

forwarding_unit FORWARDING_UNIT(
	.dREN_M(dREN_M1),
	.Equal4(\Equal4~0_combout ),
	.op_EX_1(op_EX[1]),
	.op_EX_0(op_EX[0]),
	.Equal41(\Equal4~1_combout ),
	.instruction_EX_16(instruction_EX[16]),
	.instruction_EX_17(instruction_EX[17]),
	.wsel_M_1(wsel_M[1]),
	.wsel_M_0(wsel_M[0]),
	.instruction_EX_18(instruction_EX[18]),
	.instruction_EX_19(instruction_EX[19]),
	.wsel_M_3(wsel_M[3]),
	.wsel_M_2(wsel_M[2]),
	.instruction_EX_20(instruction_EX[20]),
	.wsel_M_4(wsel_M[4]),
	.Equal0(\FORWARDING_UNIT|Equal0~2_combout ),
	.instruction_EX_22(instruction_EX[22]),
	.instruction_EX_21(instruction_EX[21]),
	.instruction_EX_24(instruction_EX[24]),
	.instruction_EX_23(instruction_EX[23]),
	.instruction_EX_25(instruction_EX[25]),
	.fuifforward_A_0(\FORWARDING_UNIT|fuif.forward_A[0]~2_combout ),
	.wsel_WB_1(wsel_WB[1]),
	.wsel_WB_0(wsel_WB[0]),
	.wsel_WB_3(wsel_WB[3]),
	.wsel_WB_2(wsel_WB[2]),
	.wsel_WB_4(wsel_WB[4]),
	.fuifforward_A_1(\FORWARDING_UNIT|fuif.forward_A[1]~5_combout ),
	.fuifbubble_lw_f(\FORWARDING_UNIT|fuif.bubble_lw_f~2_combout ),
	.regWrite_M(\regWrite_M~q ),
	.forward_B(\FORWARDING_UNIT|forward_B~0_combout ),
	.beq_EX(\beq_EX~q ),
	.bne_EX(\bne_EX~q ),
	.forward_B1(\FORWARDING_UNIT|forward_B~1_combout ),
	.Equal5(\FORWARDING_UNIT|Equal5~1_combout ),
	.regWrite_WB(\regWrite_WB~q ),
	.fuifforward_B_1(\FORWARDING_UNIT|fuif.forward_B[1]~3_combout ),
	.fuifforward_B_11(\FORWARDING_UNIT|fuif.forward_B[1]~4_combout ),
	.Equal3(\FORWARDING_UNIT|Equal3~0_combout ),
	.fuifforward_A_01(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.Equal31(\FORWARDING_UNIT|Equal3~1_combout ),
	.fuifforward_A_11(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

program_counter PROGRAM_COUNTER(
	.pc_out_3(pc_out_3),
	.pc_out_2(pc_out_2),
	.pc_out_5(pc_out_5),
	.pc_out_4(pc_out_4),
	.pc_out_7(pc_out_7),
	.pc_out_6(pc_out_6),
	.pc_out_9(pc_out_9),
	.pc_out_8(pc_out_8),
	.pc_out_11(pc_out_11),
	.pc_out_10(pc_out_10),
	.pc_out_13(pc_out_13),
	.pc_out_12(pc_out_12),
	.pc_out_15(pc_out_15),
	.pc_out_14(pc_out_14),
	.pc_out_17(pc_out_17),
	.pc_out_16(pc_out_16),
	.pc_out_19(pc_out_19),
	.pc_out_18(pc_out_18),
	.pc_out_21(pc_out_21),
	.pc_out_20(pc_out_20),
	.pc_out_23(pc_out_23),
	.pc_out_22(pc_out_22),
	.pc_out_25(pc_out_25),
	.pc_out_24(pc_out_24),
	.pc_out_27(pc_out_27),
	.pc_out_26(pc_out_26),
	.predicted_M(\predicted_M~q ),
	.pc_plus_4_2(\pc_plus_4[2]~0_combout ),
	.pc_plus_4_3(\pc_plus_4[3]~2_combout ),
	.pc_plus_4_4(\pc_plus_4[4]~4_combout ),
	.pc_plus_4_5(\pc_plus_4[5]~6_combout ),
	.pc_plus_4_6(\pc_plus_4[6]~8_combout ),
	.pc_plus_4_7(\pc_plus_4[7]~10_combout ),
	.pc_plus_4_8(\pc_plus_4[8]~12_combout ),
	.pc_plus_4_9(\pc_plus_4[9]~14_combout ),
	.pc_plus_4_10(\pc_plus_4[10]~16_combout ),
	.pc_plus_4_11(\pc_plus_4[11]~18_combout ),
	.pc_plus_4_12(\pc_plus_4[12]~20_combout ),
	.pc_plus_4_13(\pc_plus_4[13]~22_combout ),
	.pc_plus_4_14(\pc_plus_4[14]~24_combout ),
	.pc_plus_4_15(\pc_plus_4[15]~26_combout ),
	.pc_plus_4_16(\pc_plus_4[16]~28_combout ),
	.pc_plus_4_17(\pc_plus_4[17]~30_combout ),
	.pc_plus_4_18(\pc_plus_4[18]~32_combout ),
	.pc_plus_4_19(\pc_plus_4[19]~34_combout ),
	.pc_plus_4_20(\pc_plus_4[20]~36_combout ),
	.pc_plus_4_21(\pc_plus_4[21]~38_combout ),
	.pc_plus_4_22(\pc_plus_4[22]~40_combout ),
	.pc_plus_4_23(\pc_plus_4[23]~42_combout ),
	.pc_plus_4_24(\pc_plus_4[24]~44_combout ),
	.pc_plus_4_25(\pc_plus_4[25]~46_combout ),
	.pc_plus_4_26(\pc_plus_4[26]~48_combout ),
	.pc_plus_4_27(\pc_plus_4[27]~50_combout ),
	.pc_out_1(pc_out_1),
	.pc_out_0(pc_out_0),
	.pc_out_29(pc_out_29),
	.pc_out_28(pc_out_28),
	.pc_out_31(pc_out_31),
	.pc_out_30(pc_out_30),
	.j_M(\j_M~q ),
	.jal_M(\jal_M~q ),
	.branch_or_jump(\branch_or_jump~0_combout ),
	.branch_taken(\branch_taken~0_combout ),
	.jr_M(\jr_M~q ),
	.branch_or_jump1(\branch_or_jump~1_combout ),
	.predicted(\BTB|predicted~18_combout ),
	.pc_next(\pc_next~3_combout ),
	.pc_next_1(\pc_next[1]~4_combout ),
	.pc_next_0(\pc_next[0]~8_combout ),
	.pc_next_3(\pc_next[3]~10_combout ),
	.pc_next_31(\pc_next[3]~12_combout ),
	.comb(\comb~2_combout ),
	.pc_next_2(\pc_next[2]~14_combout ),
	.pc_next_21(\pc_next[2]~16_combout ),
	.pc_next_5(\pc_next[5]~18_combout ),
	.pc_next_51(\pc_next[5]~20_combout ),
	.pc_next_4(\pc_next[4]~22_combout ),
	.pc_next_41(\pc_next[4]~24_combout ),
	.pc_next_7(\pc_next[7]~26_combout ),
	.pc_next_71(\pc_next[7]~28_combout ),
	.pc_next_6(\pc_next[6]~30_combout ),
	.pc_next_61(\pc_next[6]~32_combout ),
	.pc_next_9(\pc_next[9]~34_combout ),
	.pc_next_91(\pc_next[9]~36_combout ),
	.pc_next_8(\pc_next[8]~38_combout ),
	.pc_next_81(\pc_next[8]~40_combout ),
	.pc_next_11(\pc_next[11]~42_combout ),
	.pc_next_111(\pc_next[11]~44_combout ),
	.pc_next_10(\pc_next[10]~46_combout ),
	.pc_next_101(\pc_next[10]~48_combout ),
	.pc_next_13(\pc_next[13]~50_combout ),
	.pc_next_131(\pc_next[13]~52_combout ),
	.pc_next_12(\pc_next[12]~54_combout ),
	.pc_next_121(\pc_next[12]~56_combout ),
	.pc_next_15(\pc_next[15]~58_combout ),
	.pc_next_151(\pc_next[15]~60_combout ),
	.pc_next_14(\pc_next[14]~62_combout ),
	.pc_next_141(\pc_next[14]~64_combout ),
	.pc_next_17(\pc_next[17]~66_combout ),
	.pc_next_171(\pc_next[17]~68_combout ),
	.pc_next_16(\pc_next[16]~70_combout ),
	.pc_next_161(\pc_next[16]~72_combout ),
	.pc_next_19(\pc_next[19]~74_combout ),
	.pc_next_191(\pc_next[19]~76_combout ),
	.pc_next_18(\pc_next[18]~78_combout ),
	.pc_next_181(\pc_next[18]~80_combout ),
	.pc_next_211(\pc_next[21]~82_combout ),
	.pc_next_212(\pc_next[21]~84_combout ),
	.pc_next_20(\pc_next[20]~86_combout ),
	.pc_next_201(\pc_next[20]~88_combout ),
	.pc_next_23(\pc_next[23]~90_combout ),
	.pc_next_231(\pc_next[23]~92_combout ),
	.pc_next_22(\pc_next[22]~94_combout ),
	.pc_next_221(\pc_next[22]~96_combout ),
	.pc_next_25(\pc_next[25]~98_combout ),
	.pc_next_251(\pc_next[25]~100_combout ),
	.pc_next_24(\pc_next[24]~102_combout ),
	.pc_next_241(\pc_next[24]~104_combout ),
	.pc_next_27(\pc_next[27]~106_combout ),
	.pc_next_271(\pc_next[27]~108_combout ),
	.pc_next_26(\pc_next[26]~110_combout ),
	.pc_next_261(\pc_next[26]~112_combout ),
	.pc_out_291(\PROGRAM_COUNTER|pc_out[29]~29_combout ),
	.pc_out_292(\PROGRAM_COUNTER|pc_out[29]~30_combout ),
	.pc_next_29(\pc_next[29]~117_combout ),
	.pc_next_28(\pc_next[28]~122_combout ),
	.pc_next_311(\pc_next[31]~127_combout ),
	.pc_next_30(\pc_next[30]~132_combout ),
	.comb1(\comb~3_combout ),
	.pc_out_101(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.nRST(nRST1),
	.CLK(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

control_unit CONTROL_UNIT(
	.instruction_D_31(instruction_D[31]),
	.instruction_D_28(instruction_D[28]),
	.instruction_D_30(instruction_D[30]),
	.instruction_D_29(instruction_D[29]),
	.instruction_D_27(instruction_D[27]),
	.instruction_D_26(instruction_D[26]),
	.Decoder1(\CONTROL_UNIT|Decoder1~0_combout ),
	.Decoder11(\CONTROL_UNIT|Decoder1~1_combout ),
	.Equal3(\CONTROL_UNIT|Equal3~1_combout ),
	.Equal31(\CONTROL_UNIT|Equal3~2_combout ),
	.instruction_D_5(instruction_D[5]),
	.instruction_D_0(instruction_D[0]),
	.instruction_D_3(instruction_D[3]),
	.instruction_D_2(instruction_D[2]),
	.instruction_D_1(instruction_D[1]),
	.WideOr2(\CONTROL_UNIT|WideOr2~0_combout ),
	.instruction_D_4(instruction_D[4]),
	.WideOr7(\CONTROL_UNIT|WideOr7~0_combout ),
	.WideOr6(\CONTROL_UNIT|WideOr6~0_combout ),
	.WideOr1(\CONTROL_UNIT|WideOr1~0_combout ),
	.WideOr5(\CONTROL_UNIT|WideOr5~0_combout ),
	.WideOr8(\CONTROL_UNIT|WideOr8~0_combout ),
	.WideOr4(\CONTROL_UNIT|WideOr4~0_combout ),
	.Decoder0(\CONTROL_UNIT|Decoder0~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

register_file REGISTER_FILE(
	.wsel_WB_1(wsel_WB[1]),
	.wsel_WB_0(wsel_WB[0]),
	.wsel_WB_3(wsel_WB[3]),
	.wsel_WB_2(wsel_WB[2]),
	.wsel_WB_4(wsel_WB[4]),
	.regWrite_WB(\regWrite_WB~q ),
	.wdat_WB_31(\wdat_WB[31]~3_combout ),
	.wdat_WB_30(\wdat_WB[30]~5_combout ),
	.wdat_WB_29(\wdat_WB[29]~7_combout ),
	.wdat_WB_28(\wdat_WB[28]~9_combout ),
	.wdat_WB_27(\wdat_WB[27]~11_combout ),
	.wdat_WB_26(\wdat_WB[26]~13_combout ),
	.wdat_WB_25(\wdat_WB[25]~15_combout ),
	.wdat_WB_24(\wdat_WB[24]~17_combout ),
	.wdat_WB_23(\wdat_WB[23]~19_combout ),
	.wdat_WB_22(\wdat_WB[22]~21_combout ),
	.wdat_WB_21(\wdat_WB[21]~23_combout ),
	.wdat_WB_20(\wdat_WB[20]~25_combout ),
	.wdat_WB_19(\wdat_WB[19]~27_combout ),
	.wdat_WB_18(\wdat_WB[18]~29_combout ),
	.wdat_WB_17(\wdat_WB[17]~31_combout ),
	.wdat_WB_16(\wdat_WB[16]~33_combout ),
	.wdat_WB_15(\wdat_WB[15]~35_combout ),
	.wdat_WB_14(\wdat_WB[14]~37_combout ),
	.wdat_WB_13(\wdat_WB[13]~39_combout ),
	.wdat_WB_12(\wdat_WB[12]~41_combout ),
	.wdat_WB_9(\wdat_WB[9]~43_combout ),
	.wdat_WB_8(\wdat_WB[8]~45_combout ),
	.wdat_WB_11(\wdat_WB[11]~47_combout ),
	.wdat_WB_10(\wdat_WB[10]~49_combout ),
	.wdat_WB_7(\wdat_WB[7]~51_combout ),
	.wdat_WB_6(\wdat_WB[6]~53_combout ),
	.wdat_WB_5(\wdat_WB[5]~55_combout ),
	.wdat_WB_2(\wdat_WB[2]~57_combout ),
	.wdat_WB_1(\wdat_WB[1]~59_combout ),
	.wdat_WB_0(\wdat_WB[0]~61_combout ),
	.wdat_WB_4(\wdat_WB[4]~63_combout ),
	.wdat_WB_3(\wdat_WB[3]~65_combout ),
	.instruction_D_16(instruction_D[16]),
	.instruction_D_17(instruction_D[17]),
	.instruction_D_18(instruction_D[18]),
	.instruction_D_19(instruction_D[19]),
	.instruction_D_22(instruction_D[22]),
	.instruction_D_21(instruction_D[21]),
	.instruction_D_24(instruction_D[24]),
	.instruction_D_23(instruction_D[23]),
	.Mux32(\REGISTER_FILE|Mux32~9_combout ),
	.Mux321(\REGISTER_FILE|Mux32~19_combout ),
	.Mux33(\REGISTER_FILE|Mux33~9_combout ),
	.Mux331(\REGISTER_FILE|Mux33~19_combout ),
	.Mux34(\REGISTER_FILE|Mux34~9_combout ),
	.Mux341(\REGISTER_FILE|Mux34~19_combout ),
	.Mux35(\REGISTER_FILE|Mux35~9_combout ),
	.Mux351(\REGISTER_FILE|Mux35~19_combout ),
	.Mux36(\REGISTER_FILE|Mux36~9_combout ),
	.Mux361(\REGISTER_FILE|Mux36~19_combout ),
	.Mux37(\REGISTER_FILE|Mux37~9_combout ),
	.Mux371(\REGISTER_FILE|Mux37~19_combout ),
	.Mux38(\REGISTER_FILE|Mux38~9_combout ),
	.Mux381(\REGISTER_FILE|Mux38~19_combout ),
	.Mux39(\REGISTER_FILE|Mux39~9_combout ),
	.Mux391(\REGISTER_FILE|Mux39~19_combout ),
	.Mux40(\REGISTER_FILE|Mux40~9_combout ),
	.Mux401(\REGISTER_FILE|Mux40~19_combout ),
	.Mux41(\REGISTER_FILE|Mux41~9_combout ),
	.Mux411(\REGISTER_FILE|Mux41~19_combout ),
	.Mux42(\REGISTER_FILE|Mux42~9_combout ),
	.Mux421(\REGISTER_FILE|Mux42~19_combout ),
	.Mux43(\REGISTER_FILE|Mux43~9_combout ),
	.Mux431(\REGISTER_FILE|Mux43~19_combout ),
	.Mux44(\REGISTER_FILE|Mux44~9_combout ),
	.Mux441(\REGISTER_FILE|Mux44~19_combout ),
	.Mux45(\REGISTER_FILE|Mux45~9_combout ),
	.Mux451(\REGISTER_FILE|Mux45~19_combout ),
	.Mux46(\REGISTER_FILE|Mux46~9_combout ),
	.Mux461(\REGISTER_FILE|Mux46~19_combout ),
	.Mux47(\REGISTER_FILE|Mux47~9_combout ),
	.Mux471(\REGISTER_FILE|Mux47~19_combout ),
	.Mux48(\REGISTER_FILE|Mux48~9_combout ),
	.Mux481(\REGISTER_FILE|Mux48~19_combout ),
	.Mux49(\REGISTER_FILE|Mux49~9_combout ),
	.Mux491(\REGISTER_FILE|Mux49~19_combout ),
	.Mux50(\REGISTER_FILE|Mux50~9_combout ),
	.Mux501(\REGISTER_FILE|Mux50~19_combout ),
	.Mux51(\REGISTER_FILE|Mux51~9_combout ),
	.Mux511(\REGISTER_FILE|Mux51~19_combout ),
	.Mux54(\REGISTER_FILE|Mux54~9_combout ),
	.Mux541(\REGISTER_FILE|Mux54~19_combout ),
	.Mux55(\REGISTER_FILE|Mux55~9_combout ),
	.Mux551(\REGISTER_FILE|Mux55~19_combout ),
	.Mux52(\REGISTER_FILE|Mux52~9_combout ),
	.Mux521(\REGISTER_FILE|Mux52~19_combout ),
	.Mux53(\REGISTER_FILE|Mux53~9_combout ),
	.Mux531(\REGISTER_FILE|Mux53~19_combout ),
	.Mux56(\REGISTER_FILE|Mux56~9_combout ),
	.Mux561(\REGISTER_FILE|Mux56~19_combout ),
	.Mux57(\REGISTER_FILE|Mux57~9_combout ),
	.Mux571(\REGISTER_FILE|Mux57~19_combout ),
	.Mux58(\REGISTER_FILE|Mux58~9_combout ),
	.Mux581(\REGISTER_FILE|Mux58~19_combout ),
	.Mux29(\REGISTER_FILE|Mux29~9_combout ),
	.Mux291(\REGISTER_FILE|Mux29~19_combout ),
	.Mux30(\REGISTER_FILE|Mux30~9_combout ),
	.Mux301(\REGISTER_FILE|Mux30~19_combout ),
	.Mux63(\REGISTER_FILE|Mux63~9_combout ),
	.Mux631(\REGISTER_FILE|Mux63~19_combout ),
	.Mux62(\REGISTER_FILE|Mux62~9_combout ),
	.Mux621(\REGISTER_FILE|Mux62~19_combout ),
	.Mux27(\REGISTER_FILE|Mux27~9_combout ),
	.Mux271(\REGISTER_FILE|Mux27~19_combout ),
	.Mux28(\REGISTER_FILE|Mux28~9_combout ),
	.Mux281(\REGISTER_FILE|Mux28~19_combout ),
	.Mux61(\REGISTER_FILE|Mux61~9_combout ),
	.Mux611(\REGISTER_FILE|Mux61~19_combout ),
	.Mux23(\REGISTER_FILE|Mux23~9_combout ),
	.Mux231(\REGISTER_FILE|Mux23~19_combout ),
	.Mux24(\REGISTER_FILE|Mux24~9_combout ),
	.Mux241(\REGISTER_FILE|Mux24~19_combout ),
	.Mux25(\REGISTER_FILE|Mux25~9_combout ),
	.Mux251(\REGISTER_FILE|Mux25~19_combout ),
	.Mux26(\REGISTER_FILE|Mux26~9_combout ),
	.Mux261(\REGISTER_FILE|Mux26~19_combout ),
	.Mux60(\REGISTER_FILE|Mux60~9_combout ),
	.Mux601(\REGISTER_FILE|Mux60~19_combout ),
	.Mux15(\REGISTER_FILE|Mux15~9_combout ),
	.Mux151(\REGISTER_FILE|Mux15~19_combout ),
	.Mux16(\REGISTER_FILE|Mux16~9_combout ),
	.Mux161(\REGISTER_FILE|Mux16~19_combout ),
	.Mux17(\REGISTER_FILE|Mux17~9_combout ),
	.Mux171(\REGISTER_FILE|Mux17~19_combout ),
	.Mux18(\REGISTER_FILE|Mux18~9_combout ),
	.Mux181(\REGISTER_FILE|Mux18~19_combout ),
	.Mux19(\REGISTER_FILE|Mux19~9_combout ),
	.Mux191(\REGISTER_FILE|Mux19~19_combout ),
	.Mux20(\REGISTER_FILE|Mux20~9_combout ),
	.Mux201(\REGISTER_FILE|Mux20~19_combout ),
	.Mux21(\REGISTER_FILE|Mux21~9_combout ),
	.Mux211(\REGISTER_FILE|Mux21~19_combout ),
	.Mux22(\REGISTER_FILE|Mux22~9_combout ),
	.Mux221(\REGISTER_FILE|Mux22~19_combout ),
	.Mux59(\REGISTER_FILE|Mux59~9_combout ),
	.Mux591(\REGISTER_FILE|Mux59~19_combout ),
	.Mux0(\REGISTER_FILE|Mux0~9_combout ),
	.Mux01(\REGISTER_FILE|Mux0~19_combout ),
	.Mux2(\REGISTER_FILE|Mux2~9_combout ),
	.Mux210(\REGISTER_FILE|Mux2~19_combout ),
	.Mux1(\REGISTER_FILE|Mux1~9_combout ),
	.Mux11(\REGISTER_FILE|Mux1~19_combout ),
	.Mux3(\REGISTER_FILE|Mux3~9_combout ),
	.Mux31(\REGISTER_FILE|Mux3~19_combout ),
	.Mux4(\REGISTER_FILE|Mux4~9_combout ),
	.Mux410(\REGISTER_FILE|Mux4~19_combout ),
	.Mux5(\REGISTER_FILE|Mux5~9_combout ),
	.Mux510(\REGISTER_FILE|Mux5~19_combout ),
	.Mux6(\REGISTER_FILE|Mux6~9_combout ),
	.Mux64(\REGISTER_FILE|Mux6~19_combout ),
	.Mux7(\REGISTER_FILE|Mux7~9_combout ),
	.Mux71(\REGISTER_FILE|Mux7~19_combout ),
	.Mux8(\REGISTER_FILE|Mux8~9_combout ),
	.Mux81(\REGISTER_FILE|Mux8~19_combout ),
	.Mux9(\REGISTER_FILE|Mux9~9_combout ),
	.Mux91(\REGISTER_FILE|Mux9~19_combout ),
	.Mux10(\REGISTER_FILE|Mux10~9_combout ),
	.Mux101(\REGISTER_FILE|Mux10~19_combout ),
	.Mux111(\REGISTER_FILE|Mux11~9_combout ),
	.Mux112(\REGISTER_FILE|Mux11~19_combout ),
	.Mux12(\REGISTER_FILE|Mux12~9_combout ),
	.Mux121(\REGISTER_FILE|Mux12~19_combout ),
	.Mux13(\REGISTER_FILE|Mux13~9_combout ),
	.Mux131(\REGISTER_FILE|Mux13~19_combout ),
	.Mux14(\REGISTER_FILE|Mux14~9_combout ),
	.Mux141(\REGISTER_FILE|Mux14~19_combout ),
	.Mux311(\REGISTER_FILE|Mux31~9_combout ),
	.Mux312(\REGISTER_FILE|Mux31~19_combout ),
	.nRST(nRST1),
	.CLK(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu ALU(
	.ALUOp_EX_0(ALUOp_EX[0]),
	.ALUOp_EX_1(ALUOp_EX[1]),
	.ALUOp_EX_2(ALUOp_EX[2]),
	.ALUOp_EX_3(ALUOp_EX[3]),
	.ShiftOp_EX(\ShiftOp_EX~q ),
	.portB(\portB~17_combout ),
	.portB1(\portB~20_combout ),
	.portB2(\portB~23_combout ),
	.portB3(\portB~26_combout ),
	.portB4(\portB~29_combout ),
	.portB5(\portB~32_combout ),
	.portB6(\portB~35_combout ),
	.portB7(\portB~38_combout ),
	.portB8(\portB~41_combout ),
	.portB9(\portB~44_combout ),
	.portB10(\portB~47_combout ),
	.portB11(\portB~50_combout ),
	.portB12(\portB~53_combout ),
	.portB13(\portB~56_combout ),
	.portB14(\portB~59_combout ),
	.portB15(\portB~62_combout ),
	.portB16(\portB~64_combout ),
	.portB17(\portB~66_combout ),
	.portB18(\portB~68_combout ),
	.portB19(\portB~70_combout ),
	.portB20(\portB~72_combout ),
	.portB21(\portB~73_combout ),
	.portB22(\portB~75_combout ),
	.portB23(\portB~76_combout ),
	.portB24(\portB~78_combout ),
	.portB25(\portB~80_combout ),
	.portB26(\portB~82_combout ),
	.portB27(\portB~84_combout ),
	.portB28(\portB~87_combout ),
	.fuifforward_A_1(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.portA(\portA~9_combout ),
	.portA1(\portA~12_combout ),
	.portB29(\portB~92_combout ),
	.portB30(\portB~97_combout ),
	.portA2(\portA~14_combout ),
	.wdat_WB_3(\wdat_WB[3]~65_combout ),
	.portA3(\portA~15_combout ),
	.portA4(\portA~16_combout ),
	.portB31(\portB~100_combout ),
	.portA5(\portA~17_combout ),
	.portA6(\portA~19_combout ),
	.portA7(\portA~21_combout ),
	.portA8(\portA~23_combout ),
	.portB32(\portB~103_combout ),
	.portA9(\portA~25_combout ),
	.portA10(\portA~27_combout ),
	.portA11(\portA~29_combout ),
	.portA12(\portA~31_combout ),
	.portA13(\portA~33_combout ),
	.portA14(\portA~35_combout ),
	.portA15(\portA~36_combout ),
	.portA16(\portA~37_combout ),
	.portB33(\portB~107_combout ),
	.portA17(\portA~39_combout ),
	.portA18(\portA~41_combout ),
	.portA19(\portA~43_combout ),
	.portA20(\portA~45_combout ),
	.portA21(\portA~47_combout ),
	.portA22(\portA~49_combout ),
	.portA23(\portA~51_combout ),
	.portA24(\portA~53_combout ),
	.portA25(\portA~55_combout ),
	.portA26(\portA~57_combout ),
	.portA27(\portA~59_combout ),
	.portA28(\portA~61_combout ),
	.portA29(\portA~63_combout ),
	.portA30(\portA~65_combout ),
	.portA31(\portA~67_combout ),
	.portA32(\portA~69_combout ),
	.Selector0(\ALU|Selector0~5_combout ),
	.Selector30(\ALU|Selector30~8_combout ),
	.portB34(\portB~108_combout ),
	.portB35(\portB~109_combout ),
	.Selector31(\ALU|Selector31~4_combout ),
	.Selector311(\ALU|Selector31~5_combout ),
	.Selector312(\ALU|Selector31~8_combout ),
	.Selector28(\ALU|Selector28~10_combout ),
	.Selector29(\ALU|Selector29~10_combout ),
	.Selector26(\ALU|Selector26~6_combout ),
	.Selector27(\ALU|Selector27~0_combout ),
	.Selector271(\ALU|Selector27~3_combout ),
	.Selector272(\ALU|Selector27~6_combout ),
	.Selector273(\ALU|Selector27~7_combout ),
	.Selector24(\ALU|Selector24~8_combout ),
	.Selector25(\ALU|Selector25~7_combout ),
	.Selector22(\ALU|Selector22~8_combout ),
	.Selector16(\ALU|Selector16~3_combout ),
	.Selector23(\ALU|Selector23~8_combout ),
	.Selector20(\ALU|Selector20~8_combout ),
	.Selector21(\ALU|Selector21~7_combout ),
	.Selector18(\ALU|Selector18~7_combout ),
	.Selector19(\ALU|Selector19~6_combout ),
	.ShiftLeft0(\ALU|ShiftLeft0~57_combout ),
	.Selector161(\ALU|Selector16~11_combout ),
	.Selector17(\ALU|Selector17~8_combout ),
	.Selector12(\ALU|Selector12~10_combout ),
	.Selector14(\ALU|Selector14~7_combout ),
	.Selector15(\ALU|Selector15~11_combout ),
	.Selector121(\ALU|Selector12~18_combout ),
	.Selector13(\ALU|Selector13~8_combout ),
	.Selector10(\ALU|Selector10~8_combout ),
	.Selector11(\ALU|Selector11~8_combout ),
	.Selector8(\ALU|Selector8~7_combout ),
	.Selector9(\ALU|Selector9~8_combout ),
	.Selector6(\ALU|Selector6~0_combout ),
	.Selector61(\ALU|Selector6~5_combout ),
	.Selector62(\ALU|Selector6~7_combout ),
	.Selector7(\ALU|Selector7~7_combout ),
	.Selector4(\ALU|Selector4~12_combout ),
	.Selector5(\ALU|Selector5~7_combout ),
	.Selector2(\ALU|Selector2~11_combout ),
	.Selector3(\ALU|Selector3~9_combout ),
	.Selector01(\ALU|Selector0~27_combout ),
	.Selector1(\ALU|Selector1~9_combout ),
	.Selector63(\ALU|Selector6~8_combout ),
	.Selector64(\ALU|Selector6~9_combout ),
	.Selector313(\ALU|Selector31~9_combout ),
	.Equal3(\Equal3~2_combout ),
	.ShiftRight0(\ALU|ShiftRight0~91_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X65_Y34_N31
dffeas \rdata2_EX[27] (
	.clk(CLK),
	.d(\rdata2_EX~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[27]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[27] .is_wysiwyg = "true";
defparam \rdata2_EX[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N21
dffeas \rdata2_EX[25] (
	.clk(CLK),
	.d(\rdata2_EX~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[25]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[25] .is_wysiwyg = "true";
defparam \rdata2_EX[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y34_N1
dffeas \rdata2_EX[20] (
	.clk(CLK),
	.d(\rdata2_EX~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[20]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[20] .is_wysiwyg = "true";
defparam \rdata2_EX[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N29
dffeas \rdata2_EX[13] (
	.clk(CLK),
	.d(\rdata2_EX~37_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[13]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[13] .is_wysiwyg = "true";
defparam \rdata2_EX[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N5
dffeas \rdata2_EX[8] (
	.clk(CLK),
	.d(\rdata2_EX~43_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[8]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[8] .is_wysiwyg = "true";
defparam \rdata2_EX[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N27
dffeas \rdata2_EX[11] (
	.clk(CLK),
	.d(\rdata2_EX~45_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[11]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[11] .is_wysiwyg = "true";
defparam \rdata2_EX[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N19
dffeas \rdata2_EX[10] (
	.clk(CLK),
	.d(\rdata2_EX~47_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[10]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[10] .is_wysiwyg = "true";
defparam \rdata2_EX[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N29
dffeas \rdata2_EX[7] (
	.clk(CLK),
	.d(\rdata2_EX~49_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[7]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[7] .is_wysiwyg = "true";
defparam \rdata2_EX[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N29
dffeas \rdata2_EX[5] (
	.clk(CLK),
	.d(\rdata2_EX~53_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[5]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[5] .is_wysiwyg = "true";
defparam \rdata2_EX[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N5
dffeas \rdata1_EX[2] (
	.clk(CLK),
	.d(\rdata1_EX~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[2]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[2] .is_wysiwyg = "true";
defparam \rdata1_EX[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N11
dffeas \rdata1_EX[1] (
	.clk(CLK),
	.d(\rdata1_EX~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[1]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[1] .is_wysiwyg = "true";
defparam \rdata1_EX[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N7
dffeas \rdata2_EX[0] (
	.clk(CLK),
	.d(\rdata2_EX~55_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[0]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[0] .is_wysiwyg = "true";
defparam \rdata2_EX[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N1
dffeas \rdata2_EX[1] (
	.clk(CLK),
	.d(\rdata2_EX~57_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[1]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[1] .is_wysiwyg = "true";
defparam \rdata2_EX[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N25
dffeas \rdata1_EX[4] (
	.clk(CLK),
	.d(\rdata1_EX~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[4]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[4] .is_wysiwyg = "true";
defparam \rdata1_EX[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N29
dffeas \rdata1_EX[3] (
	.clk(CLK),
	.d(\rdata1_EX~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[3]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[3] .is_wysiwyg = "true";
defparam \rdata1_EX[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N15
dffeas \rdata1_EX[8] (
	.clk(CLK),
	.d(\rdata1_EX~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[8]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[8] .is_wysiwyg = "true";
defparam \rdata1_EX[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N1
dffeas \rdata1_EX[7] (
	.clk(CLK),
	.d(\rdata1_EX~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[7]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[7] .is_wysiwyg = "true";
defparam \rdata1_EX[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N3
dffeas \rdata1_EX[6] (
	.clk(CLK),
	.d(\rdata1_EX~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[6]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[6] .is_wysiwyg = "true";
defparam \rdata1_EX[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N9
dffeas \rdata1_EX[5] (
	.clk(CLK),
	.d(\rdata1_EX~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[5]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[5] .is_wysiwyg = "true";
defparam \rdata1_EX[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N31
dffeas \rdata2_EX[3] (
	.clk(CLK),
	.d(\rdata2_EX~61_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[3]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[3] .is_wysiwyg = "true";
defparam \rdata2_EX[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N31
dffeas \rdata1_EX[16] (
	.clk(CLK),
	.d(\rdata1_EX~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[16]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[16] .is_wysiwyg = "true";
defparam \rdata1_EX[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N5
dffeas \rdata1_EX[15] (
	.clk(CLK),
	.d(\rdata1_EX~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[15]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[15] .is_wysiwyg = "true";
defparam \rdata1_EX[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N5
dffeas \rdata1_EX[14] (
	.clk(CLK),
	.d(\rdata1_EX~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[14]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[14] .is_wysiwyg = "true";
defparam \rdata1_EX[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N19
dffeas \rdata1_EX[13] (
	.clk(CLK),
	.d(\rdata1_EX~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[13]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[13] .is_wysiwyg = "true";
defparam \rdata1_EX[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N9
dffeas \rdata1_EX[12] (
	.clk(CLK),
	.d(\rdata1_EX~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[12]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[12] .is_wysiwyg = "true";
defparam \rdata1_EX[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N7
dffeas \rdata1_EX[11] (
	.clk(CLK),
	.d(\rdata1_EX~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[11]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[11] .is_wysiwyg = "true";
defparam \rdata1_EX[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y34_N3
dffeas \rdata1_EX[10] (
	.clk(CLK),
	.d(\rdata1_EX~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[10]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[10] .is_wysiwyg = "true";
defparam \rdata1_EX[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y34_N29
dffeas \rdata1_EX[9] (
	.clk(CLK),
	.d(\rdata1_EX~33_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[9]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[9] .is_wysiwyg = "true";
defparam \rdata1_EX[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y34_N15
dffeas \rdata1_EX[31] (
	.clk(CLK),
	.d(\rdata1_EX~35_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[31]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[31] .is_wysiwyg = "true";
defparam \rdata1_EX[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y34_N25
dffeas \rdata1_EX[29] (
	.clk(CLK),
	.d(\rdata1_EX~37_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[29]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[29] .is_wysiwyg = "true";
defparam \rdata1_EX[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y34_N23
dffeas \rdata1_EX[30] (
	.clk(CLK),
	.d(\rdata1_EX~39_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[30]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[30] .is_wysiwyg = "true";
defparam \rdata1_EX[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N29
dffeas \rdata1_EX[28] (
	.clk(CLK),
	.d(\rdata1_EX~41_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[28]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[28] .is_wysiwyg = "true";
defparam \rdata1_EX[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y31_N5
dffeas \rdata1_EX[27] (
	.clk(CLK),
	.d(\rdata1_EX~43_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[27]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[27] .is_wysiwyg = "true";
defparam \rdata1_EX[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y34_N21
dffeas \rdata1_EX[26] (
	.clk(CLK),
	.d(\rdata1_EX~45_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[26]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[26] .is_wysiwyg = "true";
defparam \rdata1_EX[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y31_N7
dffeas \rdata1_EX[25] (
	.clk(CLK),
	.d(\rdata1_EX~47_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[25]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[25] .is_wysiwyg = "true";
defparam \rdata1_EX[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N31
dffeas \rdata1_EX[24] (
	.clk(CLK),
	.d(\rdata1_EX~49_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[24]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[24] .is_wysiwyg = "true";
defparam \rdata1_EX[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y31_N21
dffeas \rdata1_EX[23] (
	.clk(CLK),
	.d(\rdata1_EX~51_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[23]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[23] .is_wysiwyg = "true";
defparam \rdata1_EX[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N9
dffeas \rdata1_EX[22] (
	.clk(CLK),
	.d(\rdata1_EX~53_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[22]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[22] .is_wysiwyg = "true";
defparam \rdata1_EX[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N31
dffeas \rdata1_EX[21] (
	.clk(CLK),
	.d(\rdata1_EX~55_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[21]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[21] .is_wysiwyg = "true";
defparam \rdata1_EX[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y34_N27
dffeas \rdata1_EX[20] (
	.clk(CLK),
	.d(\rdata1_EX~57_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[20]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[20] .is_wysiwyg = "true";
defparam \rdata1_EX[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N19
dffeas \rdata1_EX[19] (
	.clk(CLK),
	.d(\rdata1_EX~59_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[19]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[19] .is_wysiwyg = "true";
defparam \rdata1_EX[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y31_N3
dffeas \rdata1_EX[18] (
	.clk(CLK),
	.d(\rdata1_EX~61_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[18]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[18] .is_wysiwyg = "true";
defparam \rdata1_EX[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N13
dffeas \rdata1_EX[17] (
	.clk(CLK),
	.d(\rdata1_EX~63_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[17]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[17] .is_wysiwyg = "true";
defparam \rdata1_EX[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N13
dffeas \rdata1_M[1] (
	.clk(CLK),
	.d(\rdata1_M[1]~31_combout ),
	.asdata(\wdat_WB[1]~59_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[1]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[1] .is_wysiwyg = "true";
defparam \rdata1_M[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N23
dffeas \rdata1_M[0] (
	.clk(CLK),
	.d(\rdata1_M[0]~30_combout ),
	.asdata(\wdat_WB[0]~61_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[0]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[0] .is_wysiwyg = "true";
defparam \rdata1_M[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N29
dffeas \rdata1_M[3] (
	.clk(CLK),
	.d(\rdata1_M[3]~0_combout ),
	.asdata(\wdat_WB[3]~65_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[3]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[3] .is_wysiwyg = "true";
defparam \rdata1_M[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N2
cycloneive_lcell_comb \pc_when_branch[2]~0 (
// Equation(s):
// \pc_when_branch[2]~0_combout  = (imm_M[0] & (pc_plus_4_M[2] $ (VCC))) # (!imm_M[0] & (pc_plus_4_M[2] & VCC))
// \pc_when_branch[2]~1  = CARRY((imm_M[0] & pc_plus_4_M[2]))

	.dataa(imm_M[0]),
	.datab(pc_plus_4_M[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\pc_when_branch[2]~0_combout ),
	.cout(\pc_when_branch[2]~1 ));
// synopsys translate_off
defparam \pc_when_branch[2]~0 .lut_mask = 16'h6688;
defparam \pc_when_branch[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N4
cycloneive_lcell_comb \pc_when_branch[3]~2 (
// Equation(s):
// \pc_when_branch[3]~2_combout  = (pc_plus_4_M[3] & ((imm_M[1] & (\pc_when_branch[2]~1  & VCC)) # (!imm_M[1] & (!\pc_when_branch[2]~1 )))) # (!pc_plus_4_M[3] & ((imm_M[1] & (!\pc_when_branch[2]~1 )) # (!imm_M[1] & ((\pc_when_branch[2]~1 ) # (GND)))))
// \pc_when_branch[3]~3  = CARRY((pc_plus_4_M[3] & (!imm_M[1] & !\pc_when_branch[2]~1 )) # (!pc_plus_4_M[3] & ((!\pc_when_branch[2]~1 ) # (!imm_M[1]))))

	.dataa(pc_plus_4_M[3]),
	.datab(imm_M[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[2]~1 ),
	.combout(\pc_when_branch[3]~2_combout ),
	.cout(\pc_when_branch[3]~3 ));
// synopsys translate_off
defparam \pc_when_branch[3]~2 .lut_mask = 16'h9617;
defparam \pc_when_branch[3]~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N4
cycloneive_lcell_comb \pc_plus_4[3]~2 (
// Equation(s):
// \pc_plus_4[3]~2_combout  = (pc_out_3 & (!\pc_plus_4[2]~1 )) # (!pc_out_3 & ((\pc_plus_4[2]~1 ) # (GND)))
// \pc_plus_4[3]~3  = CARRY((!\pc_plus_4[2]~1 ) # (!pc_out_3))

	.dataa(pc_out_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[2]~1 ),
	.combout(\pc_plus_4[3]~2_combout ),
	.cout(\pc_plus_4[3]~3 ));
// synopsys translate_off
defparam \pc_plus_4[3]~2 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[3]~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X61_Y29_N25
dffeas \rdata1_M[2] (
	.clk(CLK),
	.d(\rdata1_M[2]~1_combout ),
	.asdata(\wdat_WB[2]~57_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[2]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[2] .is_wysiwyg = "true";
defparam \rdata1_M[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N6
cycloneive_lcell_comb \pc_when_branch[4]~4 (
// Equation(s):
// \pc_when_branch[4]~4_combout  = ((imm_M[2] $ (pc_plus_4_M[4] $ (!\pc_when_branch[3]~3 )))) # (GND)
// \pc_when_branch[4]~5  = CARRY((imm_M[2] & ((pc_plus_4_M[4]) # (!\pc_when_branch[3]~3 ))) # (!imm_M[2] & (pc_plus_4_M[4] & !\pc_when_branch[3]~3 )))

	.dataa(imm_M[2]),
	.datab(pc_plus_4_M[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[3]~3 ),
	.combout(\pc_when_branch[4]~4_combout ),
	.cout(\pc_when_branch[4]~5 ));
// synopsys translate_off
defparam \pc_when_branch[4]~4 .lut_mask = 16'h698E;
defparam \pc_when_branch[4]~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N8
cycloneive_lcell_comb \pc_when_branch[5]~6 (
// Equation(s):
// \pc_when_branch[5]~6_combout  = (pc_plus_4_M[5] & ((imm_M[3] & (\pc_when_branch[4]~5  & VCC)) # (!imm_M[3] & (!\pc_when_branch[4]~5 )))) # (!pc_plus_4_M[5] & ((imm_M[3] & (!\pc_when_branch[4]~5 )) # (!imm_M[3] & ((\pc_when_branch[4]~5 ) # (GND)))))
// \pc_when_branch[5]~7  = CARRY((pc_plus_4_M[5] & (!imm_M[3] & !\pc_when_branch[4]~5 )) # (!pc_plus_4_M[5] & ((!\pc_when_branch[4]~5 ) # (!imm_M[3]))))

	.dataa(pc_plus_4_M[5]),
	.datab(imm_M[3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[4]~5 ),
	.combout(\pc_when_branch[5]~6_combout ),
	.cout(\pc_when_branch[5]~7 ));
// synopsys translate_off
defparam \pc_when_branch[5]~6 .lut_mask = 16'h9617;
defparam \pc_when_branch[5]~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X62_Y28_N29
dffeas \rdata1_M[5] (
	.clk(CLK),
	.d(\rdata1_M[5]~3_combout ),
	.asdata(\wdat_WB[5]~55_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[5]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[5] .is_wysiwyg = "true";
defparam \rdata1_M[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N6
cycloneive_lcell_comb \pc_plus_4[4]~4 (
// Equation(s):
// \pc_plus_4[4]~4_combout  = (pc_out_4 & (\pc_plus_4[3]~3  $ (GND))) # (!pc_out_4 & (!\pc_plus_4[3]~3  & VCC))
// \pc_plus_4[4]~5  = CARRY((pc_out_4 & !\pc_plus_4[3]~3 ))

	.dataa(pc_out_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[3]~3 ),
	.combout(\pc_plus_4[4]~4_combout ),
	.cout(\pc_plus_4[4]~5 ));
// synopsys translate_off
defparam \pc_plus_4[4]~4 .lut_mask = 16'hA50A;
defparam \pc_plus_4[4]~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N8
cycloneive_lcell_comb \pc_plus_4[5]~6 (
// Equation(s):
// \pc_plus_4[5]~6_combout  = (pc_out_5 & (!\pc_plus_4[4]~5 )) # (!pc_out_5 & ((\pc_plus_4[4]~5 ) # (GND)))
// \pc_plus_4[5]~7  = CARRY((!\pc_plus_4[4]~5 ) # (!pc_out_5))

	.dataa(pc_out_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[4]~5 ),
	.combout(\pc_plus_4[5]~6_combout ),
	.cout(\pc_plus_4[5]~7 ));
// synopsys translate_off
defparam \pc_plus_4[5]~6 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[5]~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X62_Y28_N7
dffeas \rdata1_M[4] (
	.clk(CLK),
	.d(\rdata1_M[4]~2_combout ),
	.asdata(\wdat_WB[4]~63_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[4]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[4] .is_wysiwyg = "true";
defparam \rdata1_M[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N10
cycloneive_lcell_comb \pc_when_branch[6]~8 (
// Equation(s):
// \pc_when_branch[6]~8_combout  = ((imm_M[4] $ (pc_plus_4_M[6] $ (!\pc_when_branch[5]~7 )))) # (GND)
// \pc_when_branch[6]~9  = CARRY((imm_M[4] & ((pc_plus_4_M[6]) # (!\pc_when_branch[5]~7 ))) # (!imm_M[4] & (pc_plus_4_M[6] & !\pc_when_branch[5]~7 )))

	.dataa(imm_M[4]),
	.datab(pc_plus_4_M[6]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[5]~7 ),
	.combout(\pc_when_branch[6]~8_combout ),
	.cout(\pc_when_branch[6]~9 ));
// synopsys translate_off
defparam \pc_when_branch[6]~8 .lut_mask = 16'h698E;
defparam \pc_when_branch[6]~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N12
cycloneive_lcell_comb \pc_when_branch[7]~10 (
// Equation(s):
// \pc_when_branch[7]~10_combout  = (pc_plus_4_M[7] & ((imm_M[5] & (\pc_when_branch[6]~9  & VCC)) # (!imm_M[5] & (!\pc_when_branch[6]~9 )))) # (!pc_plus_4_M[7] & ((imm_M[5] & (!\pc_when_branch[6]~9 )) # (!imm_M[5] & ((\pc_when_branch[6]~9 ) # (GND)))))
// \pc_when_branch[7]~11  = CARRY((pc_plus_4_M[7] & (!imm_M[5] & !\pc_when_branch[6]~9 )) # (!pc_plus_4_M[7] & ((!\pc_when_branch[6]~9 ) # (!imm_M[5]))))

	.dataa(pc_plus_4_M[7]),
	.datab(imm_M[5]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[6]~9 ),
	.combout(\pc_when_branch[7]~10_combout ),
	.cout(\pc_when_branch[7]~11 ));
// synopsys translate_off
defparam \pc_when_branch[7]~10 .lut_mask = 16'h9617;
defparam \pc_when_branch[7]~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X60_Y36_N13
dffeas \rdata1_M[7] (
	.clk(CLK),
	.d(\rdata1_M[7]~5_combout ),
	.asdata(\wdat_WB[7]~51_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[7]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[7] .is_wysiwyg = "true";
defparam \rdata1_M[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N10
cycloneive_lcell_comb \pc_plus_4[6]~8 (
// Equation(s):
// \pc_plus_4[6]~8_combout  = (pc_out_6 & (\pc_plus_4[5]~7  $ (GND))) # (!pc_out_6 & (!\pc_plus_4[5]~7  & VCC))
// \pc_plus_4[6]~9  = CARRY((pc_out_6 & !\pc_plus_4[5]~7 ))

	.dataa(pc_out_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[5]~7 ),
	.combout(\pc_plus_4[6]~8_combout ),
	.cout(\pc_plus_4[6]~9 ));
// synopsys translate_off
defparam \pc_plus_4[6]~8 .lut_mask = 16'hA50A;
defparam \pc_plus_4[6]~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X65_Y35_N9
dffeas \rdata1_M[6] (
	.clk(CLK),
	.d(\rdata1_M[6]~4_combout ),
	.asdata(\wdat_WB[6]~53_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[6]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[6] .is_wysiwyg = "true";
defparam \rdata1_M[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N14
cycloneive_lcell_comb \pc_when_branch[8]~12 (
// Equation(s):
// \pc_when_branch[8]~12_combout  = ((imm_M[6] $ (pc_plus_4_M[8] $ (!\pc_when_branch[7]~11 )))) # (GND)
// \pc_when_branch[8]~13  = CARRY((imm_M[6] & ((pc_plus_4_M[8]) # (!\pc_when_branch[7]~11 ))) # (!imm_M[6] & (pc_plus_4_M[8] & !\pc_when_branch[7]~11 )))

	.dataa(imm_M[6]),
	.datab(pc_plus_4_M[8]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[7]~11 ),
	.combout(\pc_when_branch[8]~12_combout ),
	.cout(\pc_when_branch[8]~13 ));
// synopsys translate_off
defparam \pc_when_branch[8]~12 .lut_mask = 16'h698E;
defparam \pc_when_branch[8]~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N16
cycloneive_lcell_comb \pc_when_branch[9]~14 (
// Equation(s):
// \pc_when_branch[9]~14_combout  = (imm_M[7] & ((pc_plus_4_M[9] & (\pc_when_branch[8]~13  & VCC)) # (!pc_plus_4_M[9] & (!\pc_when_branch[8]~13 )))) # (!imm_M[7] & ((pc_plus_4_M[9] & (!\pc_when_branch[8]~13 )) # (!pc_plus_4_M[9] & ((\pc_when_branch[8]~13 ) # 
// (GND)))))
// \pc_when_branch[9]~15  = CARRY((imm_M[7] & (!pc_plus_4_M[9] & !\pc_when_branch[8]~13 )) # (!imm_M[7] & ((!\pc_when_branch[8]~13 ) # (!pc_plus_4_M[9]))))

	.dataa(imm_M[7]),
	.datab(pc_plus_4_M[9]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[8]~13 ),
	.combout(\pc_when_branch[9]~14_combout ),
	.cout(\pc_when_branch[9]~15 ));
// synopsys translate_off
defparam \pc_when_branch[9]~14 .lut_mask = 16'h9617;
defparam \pc_when_branch[9]~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X60_Y36_N3
dffeas \rdata1_M[9] (
	.clk(CLK),
	.d(\rdata1_M[9]~7_combout ),
	.asdata(\wdat_WB[9]~43_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[9]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[9] .is_wysiwyg = "true";
defparam \rdata1_M[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N14
cycloneive_lcell_comb \pc_plus_4[8]~12 (
// Equation(s):
// \pc_plus_4[8]~12_combout  = (pc_out_8 & (\pc_plus_4[7]~11  $ (GND))) # (!pc_out_8 & (!\pc_plus_4[7]~11  & VCC))
// \pc_plus_4[8]~13  = CARRY((pc_out_8 & !\pc_plus_4[7]~11 ))

	.dataa(pc_out_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[7]~11 ),
	.combout(\pc_plus_4[8]~12_combout ),
	.cout(\pc_plus_4[8]~13 ));
// synopsys translate_off
defparam \pc_plus_4[8]~12 .lut_mask = 16'hA50A;
defparam \pc_plus_4[8]~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N16
cycloneive_lcell_comb \pc_plus_4[9]~14 (
// Equation(s):
// \pc_plus_4[9]~14_combout  = (pc_out_9 & (!\pc_plus_4[8]~13 )) # (!pc_out_9 & ((\pc_plus_4[8]~13 ) # (GND)))
// \pc_plus_4[9]~15  = CARRY((!\pc_plus_4[8]~13 ) # (!pc_out_9))

	.dataa(pc_out_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[8]~13 ),
	.combout(\pc_plus_4[9]~14_combout ),
	.cout(\pc_plus_4[9]~15 ));
// synopsys translate_off
defparam \pc_plus_4[9]~14 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[9]~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X60_Y36_N25
dffeas \rdata1_M[8] (
	.clk(CLK),
	.d(\rdata1_M[8]~6_combout ),
	.asdata(\wdat_WB[8]~45_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[8]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[8] .is_wysiwyg = "true";
defparam \rdata1_M[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N18
cycloneive_lcell_comb \pc_when_branch[10]~16 (
// Equation(s):
// \pc_when_branch[10]~16_combout  = ((pc_plus_4_M[10] $ (imm_M[8] $ (!\pc_when_branch[9]~15 )))) # (GND)
// \pc_when_branch[10]~17  = CARRY((pc_plus_4_M[10] & ((imm_M[8]) # (!\pc_when_branch[9]~15 ))) # (!pc_plus_4_M[10] & (imm_M[8] & !\pc_when_branch[9]~15 )))

	.dataa(pc_plus_4_M[10]),
	.datab(imm_M[8]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[9]~15 ),
	.combout(\pc_when_branch[10]~16_combout ),
	.cout(\pc_when_branch[10]~17 ));
// synopsys translate_off
defparam \pc_when_branch[10]~16 .lut_mask = 16'h698E;
defparam \pc_when_branch[10]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N20
cycloneive_lcell_comb \pc_when_branch[11]~18 (
// Equation(s):
// \pc_when_branch[11]~18_combout  = (pc_plus_4_M[11] & ((imm_M[9] & (\pc_when_branch[10]~17  & VCC)) # (!imm_M[9] & (!\pc_when_branch[10]~17 )))) # (!pc_plus_4_M[11] & ((imm_M[9] & (!\pc_when_branch[10]~17 )) # (!imm_M[9] & ((\pc_when_branch[10]~17 ) # 
// (GND)))))
// \pc_when_branch[11]~19  = CARRY((pc_plus_4_M[11] & (!imm_M[9] & !\pc_when_branch[10]~17 )) # (!pc_plus_4_M[11] & ((!\pc_when_branch[10]~17 ) # (!imm_M[9]))))

	.dataa(pc_plus_4_M[11]),
	.datab(imm_M[9]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[10]~17 ),
	.combout(\pc_when_branch[11]~18_combout ),
	.cout(\pc_when_branch[11]~19 ));
// synopsys translate_off
defparam \pc_when_branch[11]~18 .lut_mask = 16'h9617;
defparam \pc_when_branch[11]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X62_Y28_N1
dffeas \rdata1_M[11] (
	.clk(CLK),
	.d(\rdata1_M[11]~9_combout ),
	.asdata(\wdat_WB[11]~47_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[11]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[11] .is_wysiwyg = "true";
defparam \rdata1_M[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N18
cycloneive_lcell_comb \pc_plus_4[10]~16 (
// Equation(s):
// \pc_plus_4[10]~16_combout  = (pc_out_10 & (\pc_plus_4[9]~15  $ (GND))) # (!pc_out_10 & (!\pc_plus_4[9]~15  & VCC))
// \pc_plus_4[10]~17  = CARRY((pc_out_10 & !\pc_plus_4[9]~15 ))

	.dataa(pc_out_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[9]~15 ),
	.combout(\pc_plus_4[10]~16_combout ),
	.cout(\pc_plus_4[10]~17 ));
// synopsys translate_off
defparam \pc_plus_4[10]~16 .lut_mask = 16'hA50A;
defparam \pc_plus_4[10]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N20
cycloneive_lcell_comb \pc_plus_4[11]~18 (
// Equation(s):
// \pc_plus_4[11]~18_combout  = (pc_out_11 & (!\pc_plus_4[10]~17 )) # (!pc_out_11 & ((\pc_plus_4[10]~17 ) # (GND)))
// \pc_plus_4[11]~19  = CARRY((!\pc_plus_4[10]~17 ) # (!pc_out_11))

	.dataa(pc_out_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[10]~17 ),
	.combout(\pc_plus_4[11]~18_combout ),
	.cout(\pc_plus_4[11]~19 ));
// synopsys translate_off
defparam \pc_plus_4[11]~18 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[11]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X61_Y34_N13
dffeas \rdata1_M[10] (
	.clk(CLK),
	.d(\rdata1_M[10]~8_combout ),
	.asdata(\wdat_WB[10]~49_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[10]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[10] .is_wysiwyg = "true";
defparam \rdata1_M[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N22
cycloneive_lcell_comb \pc_when_branch[12]~20 (
// Equation(s):
// \pc_when_branch[12]~20_combout  = ((pc_plus_4_M[12] $ (imm_M[10] $ (!\pc_when_branch[11]~19 )))) # (GND)
// \pc_when_branch[12]~21  = CARRY((pc_plus_4_M[12] & ((imm_M[10]) # (!\pc_when_branch[11]~19 ))) # (!pc_plus_4_M[12] & (imm_M[10] & !\pc_when_branch[11]~19 )))

	.dataa(pc_plus_4_M[12]),
	.datab(imm_M[10]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[11]~19 ),
	.combout(\pc_when_branch[12]~20_combout ),
	.cout(\pc_when_branch[12]~21 ));
// synopsys translate_off
defparam \pc_when_branch[12]~20 .lut_mask = 16'h698E;
defparam \pc_when_branch[12]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N24
cycloneive_lcell_comb \pc_when_branch[13]~22 (
// Equation(s):
// \pc_when_branch[13]~22_combout  = (pc_plus_4_M[13] & ((imm_M[11] & (\pc_when_branch[12]~21  & VCC)) # (!imm_M[11] & (!\pc_when_branch[12]~21 )))) # (!pc_plus_4_M[13] & ((imm_M[11] & (!\pc_when_branch[12]~21 )) # (!imm_M[11] & ((\pc_when_branch[12]~21 ) # 
// (GND)))))
// \pc_when_branch[13]~23  = CARRY((pc_plus_4_M[13] & (!imm_M[11] & !\pc_when_branch[12]~21 )) # (!pc_plus_4_M[13] & ((!\pc_when_branch[12]~21 ) # (!imm_M[11]))))

	.dataa(pc_plus_4_M[13]),
	.datab(imm_M[11]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[12]~21 ),
	.combout(\pc_when_branch[13]~22_combout ),
	.cout(\pc_when_branch[13]~23 ));
// synopsys translate_off
defparam \pc_when_branch[13]~22 .lut_mask = 16'h9617;
defparam \pc_when_branch[13]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X59_Y35_N5
dffeas \rdata1_M[13] (
	.clk(CLK),
	.d(\rdata1_M[13]~11_combout ),
	.asdata(\wdat_WB[13]~39_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[13]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[13] .is_wysiwyg = "true";
defparam \rdata1_M[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N22
cycloneive_lcell_comb \pc_plus_4[12]~20 (
// Equation(s):
// \pc_plus_4[12]~20_combout  = (pc_out_12 & (\pc_plus_4[11]~19  $ (GND))) # (!pc_out_12 & (!\pc_plus_4[11]~19  & VCC))
// \pc_plus_4[12]~21  = CARRY((pc_out_12 & !\pc_plus_4[11]~19 ))

	.dataa(gnd),
	.datab(pc_out_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[11]~19 ),
	.combout(\pc_plus_4[12]~20_combout ),
	.cout(\pc_plus_4[12]~21 ));
// synopsys translate_off
defparam \pc_plus_4[12]~20 .lut_mask = 16'hC30C;
defparam \pc_plus_4[12]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N24
cycloneive_lcell_comb \pc_plus_4[13]~22 (
// Equation(s):
// \pc_plus_4[13]~22_combout  = (pc_out_13 & (!\pc_plus_4[12]~21 )) # (!pc_out_13 & ((\pc_plus_4[12]~21 ) # (GND)))
// \pc_plus_4[13]~23  = CARRY((!\pc_plus_4[12]~21 ) # (!pc_out_13))

	.dataa(pc_out_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[12]~21 ),
	.combout(\pc_plus_4[13]~22_combout ),
	.cout(\pc_plus_4[13]~23 ));
// synopsys translate_off
defparam \pc_plus_4[13]~22 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[13]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X59_Y37_N29
dffeas \rdata1_M[12] (
	.clk(CLK),
	.d(\rdata1_M[12]~10_combout ),
	.asdata(\wdat_WB[12]~41_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[12]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[12] .is_wysiwyg = "true";
defparam \rdata1_M[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N26
cycloneive_lcell_comb \pc_when_branch[14]~24 (
// Equation(s):
// \pc_when_branch[14]~24_combout  = ((imm_M[12] $ (pc_plus_4_M[14] $ (!\pc_when_branch[13]~23 )))) # (GND)
// \pc_when_branch[14]~25  = CARRY((imm_M[12] & ((pc_plus_4_M[14]) # (!\pc_when_branch[13]~23 ))) # (!imm_M[12] & (pc_plus_4_M[14] & !\pc_when_branch[13]~23 )))

	.dataa(imm_M[12]),
	.datab(pc_plus_4_M[14]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[13]~23 ),
	.combout(\pc_when_branch[14]~24_combout ),
	.cout(\pc_when_branch[14]~25 ));
// synopsys translate_off
defparam \pc_when_branch[14]~24 .lut_mask = 16'h698E;
defparam \pc_when_branch[14]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N28
cycloneive_lcell_comb \pc_when_branch[15]~26 (
// Equation(s):
// \pc_when_branch[15]~26_combout  = (pc_plus_4_M[15] & ((imm_M[13] & (\pc_when_branch[14]~25  & VCC)) # (!imm_M[13] & (!\pc_when_branch[14]~25 )))) # (!pc_plus_4_M[15] & ((imm_M[13] & (!\pc_when_branch[14]~25 )) # (!imm_M[13] & ((\pc_when_branch[14]~25 ) # 
// (GND)))))
// \pc_when_branch[15]~27  = CARRY((pc_plus_4_M[15] & (!imm_M[13] & !\pc_when_branch[14]~25 )) # (!pc_plus_4_M[15] & ((!\pc_when_branch[14]~25 ) # (!imm_M[13]))))

	.dataa(pc_plus_4_M[15]),
	.datab(imm_M[13]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[14]~25 ),
	.combout(\pc_when_branch[15]~26_combout ),
	.cout(\pc_when_branch[15]~27 ));
// synopsys translate_off
defparam \pc_when_branch[15]~26 .lut_mask = 16'h9617;
defparam \pc_when_branch[15]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X62_Y28_N27
dffeas \rdata1_M[15] (
	.clk(CLK),
	.d(\rdata1_M[15]~13_combout ),
	.asdata(\wdat_WB[15]~35_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[15]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[15] .is_wysiwyg = "true";
defparam \rdata1_M[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N26
cycloneive_lcell_comb \pc_plus_4[14]~24 (
// Equation(s):
// \pc_plus_4[14]~24_combout  = (pc_out_14 & (\pc_plus_4[13]~23  $ (GND))) # (!pc_out_14 & (!\pc_plus_4[13]~23  & VCC))
// \pc_plus_4[14]~25  = CARRY((pc_out_14 & !\pc_plus_4[13]~23 ))

	.dataa(pc_out_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[13]~23 ),
	.combout(\pc_plus_4[14]~24_combout ),
	.cout(\pc_plus_4[14]~25 ));
// synopsys translate_off
defparam \pc_plus_4[14]~24 .lut_mask = 16'hA50A;
defparam \pc_plus_4[14]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N28
cycloneive_lcell_comb \pc_plus_4[15]~26 (
// Equation(s):
// \pc_plus_4[15]~26_combout  = (pc_out_15 & (!\pc_plus_4[14]~25 )) # (!pc_out_15 & ((\pc_plus_4[14]~25 ) # (GND)))
// \pc_plus_4[15]~27  = CARRY((!\pc_plus_4[14]~25 ) # (!pc_out_15))

	.dataa(gnd),
	.datab(pc_out_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[14]~25 ),
	.combout(\pc_plus_4[15]~26_combout ),
	.cout(\pc_plus_4[15]~27 ));
// synopsys translate_off
defparam \pc_plus_4[15]~26 .lut_mask = 16'h3C3F;
defparam \pc_plus_4[15]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X62_Y28_N17
dffeas \rdata1_M[14] (
	.clk(CLK),
	.d(\rdata1_M[14]~12_combout ),
	.asdata(\wdat_WB[14]~37_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[14]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[14] .is_wysiwyg = "true";
defparam \rdata1_M[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N30
cycloneive_lcell_comb \pc_when_branch[16]~28 (
// Equation(s):
// \pc_when_branch[16]~28_combout  = ((imm_M[14] $ (pc_plus_4_M[16] $ (!\pc_when_branch[15]~27 )))) # (GND)
// \pc_when_branch[16]~29  = CARRY((imm_M[14] & ((pc_plus_4_M[16]) # (!\pc_when_branch[15]~27 ))) # (!imm_M[14] & (pc_plus_4_M[16] & !\pc_when_branch[15]~27 )))

	.dataa(imm_M[14]),
	.datab(pc_plus_4_M[16]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[15]~27 ),
	.combout(\pc_when_branch[16]~28_combout ),
	.cout(\pc_when_branch[16]~29 ));
// synopsys translate_off
defparam \pc_when_branch[16]~28 .lut_mask = 16'h698E;
defparam \pc_when_branch[16]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N0
cycloneive_lcell_comb \pc_when_branch[17]~30 (
// Equation(s):
// \pc_when_branch[17]~30_combout  = (imm_M[15] & ((pc_plus_4_M[17] & (\pc_when_branch[16]~29  & VCC)) # (!pc_plus_4_M[17] & (!\pc_when_branch[16]~29 )))) # (!imm_M[15] & ((pc_plus_4_M[17] & (!\pc_when_branch[16]~29 )) # (!pc_plus_4_M[17] & 
// ((\pc_when_branch[16]~29 ) # (GND)))))
// \pc_when_branch[17]~31  = CARRY((imm_M[15] & (!pc_plus_4_M[17] & !\pc_when_branch[16]~29 )) # (!imm_M[15] & ((!\pc_when_branch[16]~29 ) # (!pc_plus_4_M[17]))))

	.dataa(imm_M[15]),
	.datab(pc_plus_4_M[17]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[16]~29 ),
	.combout(\pc_when_branch[17]~30_combout ),
	.cout(\pc_when_branch[17]~31 ));
// synopsys translate_off
defparam \pc_when_branch[17]~30 .lut_mask = 16'h9617;
defparam \pc_when_branch[17]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X62_Y28_N3
dffeas \rdata1_M[17] (
	.clk(CLK),
	.d(\rdata1_M[17]~15_combout ),
	.asdata(\wdat_WB[17]~31_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[17]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[17] .is_wysiwyg = "true";
defparam \rdata1_M[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N30
cycloneive_lcell_comb \pc_plus_4[16]~28 (
// Equation(s):
// \pc_plus_4[16]~28_combout  = (pc_out_16 & (\pc_plus_4[15]~27  $ (GND))) # (!pc_out_16 & (!\pc_plus_4[15]~27  & VCC))
// \pc_plus_4[16]~29  = CARRY((pc_out_16 & !\pc_plus_4[15]~27 ))

	.dataa(pc_out_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[15]~27 ),
	.combout(\pc_plus_4[16]~28_combout ),
	.cout(\pc_plus_4[16]~29 ));
// synopsys translate_off
defparam \pc_plus_4[16]~28 .lut_mask = 16'hA50A;
defparam \pc_plus_4[16]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X60_Y37_N23
dffeas \rdata1_M[16] (
	.clk(CLK),
	.d(\rdata1_M[16]~14_combout ),
	.asdata(\wdat_WB[16]~33_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[16]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[16] .is_wysiwyg = "true";
defparam \rdata1_M[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N2
cycloneive_lcell_comb \pc_when_branch[18]~32 (
// Equation(s):
// \pc_when_branch[18]~32_combout  = ((imm_M[15] $ (pc_plus_4_M[18] $ (!\pc_when_branch[17]~31 )))) # (GND)
// \pc_when_branch[18]~33  = CARRY((imm_M[15] & ((pc_plus_4_M[18]) # (!\pc_when_branch[17]~31 ))) # (!imm_M[15] & (pc_plus_4_M[18] & !\pc_when_branch[17]~31 )))

	.dataa(imm_M[15]),
	.datab(pc_plus_4_M[18]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[17]~31 ),
	.combout(\pc_when_branch[18]~32_combout ),
	.cout(\pc_when_branch[18]~33 ));
// synopsys translate_off
defparam \pc_when_branch[18]~32 .lut_mask = 16'h698E;
defparam \pc_when_branch[18]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N4
cycloneive_lcell_comb \pc_when_branch[19]~34 (
// Equation(s):
// \pc_when_branch[19]~34_combout  = (imm_M[15] & ((pc_plus_4_M[19] & (\pc_when_branch[18]~33  & VCC)) # (!pc_plus_4_M[19] & (!\pc_when_branch[18]~33 )))) # (!imm_M[15] & ((pc_plus_4_M[19] & (!\pc_when_branch[18]~33 )) # (!pc_plus_4_M[19] & 
// ((\pc_when_branch[18]~33 ) # (GND)))))
// \pc_when_branch[19]~35  = CARRY((imm_M[15] & (!pc_plus_4_M[19] & !\pc_when_branch[18]~33 )) # (!imm_M[15] & ((!\pc_when_branch[18]~33 ) # (!pc_plus_4_M[19]))))

	.dataa(imm_M[15]),
	.datab(pc_plus_4_M[19]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[18]~33 ),
	.combout(\pc_when_branch[19]~34_combout ),
	.cout(\pc_when_branch[19]~35 ));
// synopsys translate_off
defparam \pc_when_branch[19]~34 .lut_mask = 16'h9617;
defparam \pc_when_branch[19]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X59_Y37_N11
dffeas \rdata1_M[19] (
	.clk(CLK),
	.d(\rdata1_M[19]~17_combout ),
	.asdata(\wdat_WB[19]~27_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[19]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[19] .is_wysiwyg = "true";
defparam \rdata1_M[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N2
cycloneive_lcell_comb \pc_plus_4[18]~32 (
// Equation(s):
// \pc_plus_4[18]~32_combout  = (pc_out_18 & (\pc_plus_4[17]~31  $ (GND))) # (!pc_out_18 & (!\pc_plus_4[17]~31  & VCC))
// \pc_plus_4[18]~33  = CARRY((pc_out_18 & !\pc_plus_4[17]~31 ))

	.dataa(gnd),
	.datab(pc_out_18),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[17]~31 ),
	.combout(\pc_plus_4[18]~32_combout ),
	.cout(\pc_plus_4[18]~33 ));
// synopsys translate_off
defparam \pc_plus_4[18]~32 .lut_mask = 16'hC30C;
defparam \pc_plus_4[18]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X59_Y38_N1
dffeas \rdata1_M[18] (
	.clk(CLK),
	.d(\rdata1_M[18]~16_combout ),
	.asdata(\wdat_WB[18]~29_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[18]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[18] .is_wysiwyg = "true";
defparam \rdata1_M[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N6
cycloneive_lcell_comb \pc_when_branch[20]~36 (
// Equation(s):
// \pc_when_branch[20]~36_combout  = ((imm_M[15] $ (pc_plus_4_M[20] $ (!\pc_when_branch[19]~35 )))) # (GND)
// \pc_when_branch[20]~37  = CARRY((imm_M[15] & ((pc_plus_4_M[20]) # (!\pc_when_branch[19]~35 ))) # (!imm_M[15] & (pc_plus_4_M[20] & !\pc_when_branch[19]~35 )))

	.dataa(imm_M[15]),
	.datab(pc_plus_4_M[20]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[19]~35 ),
	.combout(\pc_when_branch[20]~36_combout ),
	.cout(\pc_when_branch[20]~37 ));
// synopsys translate_off
defparam \pc_when_branch[20]~36 .lut_mask = 16'h698E;
defparam \pc_when_branch[20]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N8
cycloneive_lcell_comb \pc_when_branch[21]~38 (
// Equation(s):
// \pc_when_branch[21]~38_combout  = (imm_M[15] & ((pc_plus_4_M[21] & (\pc_when_branch[20]~37  & VCC)) # (!pc_plus_4_M[21] & (!\pc_when_branch[20]~37 )))) # (!imm_M[15] & ((pc_plus_4_M[21] & (!\pc_when_branch[20]~37 )) # (!pc_plus_4_M[21] & 
// ((\pc_when_branch[20]~37 ) # (GND)))))
// \pc_when_branch[21]~39  = CARRY((imm_M[15] & (!pc_plus_4_M[21] & !\pc_when_branch[20]~37 )) # (!imm_M[15] & ((!\pc_when_branch[20]~37 ) # (!pc_plus_4_M[21]))))

	.dataa(imm_M[15]),
	.datab(pc_plus_4_M[21]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[20]~37 ),
	.combout(\pc_when_branch[21]~38_combout ),
	.cout(\pc_when_branch[21]~39 ));
// synopsys translate_off
defparam \pc_when_branch[21]~38 .lut_mask = 16'h9617;
defparam \pc_when_branch[21]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X61_Y29_N27
dffeas \rdata1_M[21] (
	.clk(CLK),
	.d(\rdata1_M[21]~19_combout ),
	.asdata(\wdat_WB[21]~23_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[21]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[21] .is_wysiwyg = "true";
defparam \rdata1_M[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N8
cycloneive_lcell_comb \pc_plus_4[21]~38 (
// Equation(s):
// \pc_plus_4[21]~38_combout  = (pc_out_21 & (!\pc_plus_4[20]~37 )) # (!pc_out_21 & ((\pc_plus_4[20]~37 ) # (GND)))
// \pc_plus_4[21]~39  = CARRY((!\pc_plus_4[20]~37 ) # (!pc_out_21))

	.dataa(pc_out_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[20]~37 ),
	.combout(\pc_plus_4[21]~38_combout ),
	.cout(\pc_plus_4[21]~39 ));
// synopsys translate_off
defparam \pc_plus_4[21]~38 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[21]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X59_Y37_N9
dffeas \rdata1_M[20] (
	.clk(CLK),
	.d(\rdata1_M[20]~18_combout ),
	.asdata(\wdat_WB[20]~25_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[20]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[20] .is_wysiwyg = "true";
defparam \rdata1_M[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N10
cycloneive_lcell_comb \pc_when_branch[22]~40 (
// Equation(s):
// \pc_when_branch[22]~40_combout  = ((imm_M[15] $ (pc_plus_4_M[22] $ (!\pc_when_branch[21]~39 )))) # (GND)
// \pc_when_branch[22]~41  = CARRY((imm_M[15] & ((pc_plus_4_M[22]) # (!\pc_when_branch[21]~39 ))) # (!imm_M[15] & (pc_plus_4_M[22] & !\pc_when_branch[21]~39 )))

	.dataa(imm_M[15]),
	.datab(pc_plus_4_M[22]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[21]~39 ),
	.combout(\pc_when_branch[22]~40_combout ),
	.cout(\pc_when_branch[22]~41 ));
// synopsys translate_off
defparam \pc_when_branch[22]~40 .lut_mask = 16'h698E;
defparam \pc_when_branch[22]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N12
cycloneive_lcell_comb \pc_when_branch[23]~42 (
// Equation(s):
// \pc_when_branch[23]~42_combout  = (imm_M[15] & ((pc_plus_4_M[23] & (\pc_when_branch[22]~41  & VCC)) # (!pc_plus_4_M[23] & (!\pc_when_branch[22]~41 )))) # (!imm_M[15] & ((pc_plus_4_M[23] & (!\pc_when_branch[22]~41 )) # (!pc_plus_4_M[23] & 
// ((\pc_when_branch[22]~41 ) # (GND)))))
// \pc_when_branch[23]~43  = CARRY((imm_M[15] & (!pc_plus_4_M[23] & !\pc_when_branch[22]~41 )) # (!imm_M[15] & ((!\pc_when_branch[22]~41 ) # (!pc_plus_4_M[23]))))

	.dataa(imm_M[15]),
	.datab(pc_plus_4_M[23]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[22]~41 ),
	.combout(\pc_when_branch[23]~42_combout ),
	.cout(\pc_when_branch[23]~43 ));
// synopsys translate_off
defparam \pc_when_branch[23]~42 .lut_mask = 16'h9617;
defparam \pc_when_branch[23]~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X62_Y28_N25
dffeas \rdata1_M[23] (
	.clk(CLK),
	.d(\rdata1_M[23]~21_combout ),
	.asdata(\wdat_WB[23]~19_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[23]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[23] .is_wysiwyg = "true";
defparam \rdata1_M[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N10
cycloneive_lcell_comb \pc_plus_4[22]~40 (
// Equation(s):
// \pc_plus_4[22]~40_combout  = (pc_out_22 & (\pc_plus_4[21]~39  $ (GND))) # (!pc_out_22 & (!\pc_plus_4[21]~39  & VCC))
// \pc_plus_4[22]~41  = CARRY((pc_out_22 & !\pc_plus_4[21]~39 ))

	.dataa(pc_out_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[21]~39 ),
	.combout(\pc_plus_4[22]~40_combout ),
	.cout(\pc_plus_4[22]~41 ));
// synopsys translate_off
defparam \pc_plus_4[22]~40 .lut_mask = 16'hA50A;
defparam \pc_plus_4[22]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X59_Y35_N11
dffeas \rdata1_M[22] (
	.clk(CLK),
	.d(\rdata1_M[22]~20_combout ),
	.asdata(\wdat_WB[22]~21_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[22]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[22] .is_wysiwyg = "true";
defparam \rdata1_M[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N14
cycloneive_lcell_comb \pc_when_branch[24]~44 (
// Equation(s):
// \pc_when_branch[24]~44_combout  = ((pc_plus_4_M[24] $ (imm_M[15] $ (!\pc_when_branch[23]~43 )))) # (GND)
// \pc_when_branch[24]~45  = CARRY((pc_plus_4_M[24] & ((imm_M[15]) # (!\pc_when_branch[23]~43 ))) # (!pc_plus_4_M[24] & (imm_M[15] & !\pc_when_branch[23]~43 )))

	.dataa(pc_plus_4_M[24]),
	.datab(imm_M[15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[23]~43 ),
	.combout(\pc_when_branch[24]~44_combout ),
	.cout(\pc_when_branch[24]~45 ));
// synopsys translate_off
defparam \pc_when_branch[24]~44 .lut_mask = 16'h698E;
defparam \pc_when_branch[24]~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N16
cycloneive_lcell_comb \pc_when_branch[25]~46 (
// Equation(s):
// \pc_when_branch[25]~46_combout  = (pc_plus_4_M[25] & ((imm_M[15] & (\pc_when_branch[24]~45  & VCC)) # (!imm_M[15] & (!\pc_when_branch[24]~45 )))) # (!pc_plus_4_M[25] & ((imm_M[15] & (!\pc_when_branch[24]~45 )) # (!imm_M[15] & ((\pc_when_branch[24]~45 ) # 
// (GND)))))
// \pc_when_branch[25]~47  = CARRY((pc_plus_4_M[25] & (!imm_M[15] & !\pc_when_branch[24]~45 )) # (!pc_plus_4_M[25] & ((!\pc_when_branch[24]~45 ) # (!imm_M[15]))))

	.dataa(pc_plus_4_M[25]),
	.datab(imm_M[15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[24]~45 ),
	.combout(\pc_when_branch[25]~46_combout ),
	.cout(\pc_when_branch[25]~47 ));
// synopsys translate_off
defparam \pc_when_branch[25]~46 .lut_mask = 16'h9617;
defparam \pc_when_branch[25]~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X60_Y37_N1
dffeas \rdata1_M[25] (
	.clk(CLK),
	.d(\rdata1_M[25]~23_combout ),
	.asdata(\wdat_WB[25]~15_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[25]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[25] .is_wysiwyg = "true";
defparam \rdata1_M[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N14
cycloneive_lcell_comb \pc_plus_4[24]~44 (
// Equation(s):
// \pc_plus_4[24]~44_combout  = (pc_out_24 & (\pc_plus_4[23]~43  $ (GND))) # (!pc_out_24 & (!\pc_plus_4[23]~43  & VCC))
// \pc_plus_4[24]~45  = CARRY((pc_out_24 & !\pc_plus_4[23]~43 ))

	.dataa(gnd),
	.datab(pc_out_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[23]~43 ),
	.combout(\pc_plus_4[24]~44_combout ),
	.cout(\pc_plus_4[24]~45 ));
// synopsys translate_off
defparam \pc_plus_4[24]~44 .lut_mask = 16'hC30C;
defparam \pc_plus_4[24]~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X59_Y32_N13
dffeas \rdata1_M[24] (
	.clk(CLK),
	.d(\rdata1_M[24]~22_combout ),
	.asdata(\wdat_WB[24]~17_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[24]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[24] .is_wysiwyg = "true";
defparam \rdata1_M[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N18
cycloneive_lcell_comb \pc_when_branch[26]~48 (
// Equation(s):
// \pc_when_branch[26]~48_combout  = ((pc_plus_4_M[26] $ (imm_M[15] $ (!\pc_when_branch[25]~47 )))) # (GND)
// \pc_when_branch[26]~49  = CARRY((pc_plus_4_M[26] & ((imm_M[15]) # (!\pc_when_branch[25]~47 ))) # (!pc_plus_4_M[26] & (imm_M[15] & !\pc_when_branch[25]~47 )))

	.dataa(pc_plus_4_M[26]),
	.datab(imm_M[15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[25]~47 ),
	.combout(\pc_when_branch[26]~48_combout ),
	.cout(\pc_when_branch[26]~49 ));
// synopsys translate_off
defparam \pc_when_branch[26]~48 .lut_mask = 16'h698E;
defparam \pc_when_branch[26]~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N20
cycloneive_lcell_comb \pc_when_branch[27]~50 (
// Equation(s):
// \pc_when_branch[27]~50_combout  = (pc_plus_4_M[27] & ((imm_M[15] & (\pc_when_branch[26]~49  & VCC)) # (!imm_M[15] & (!\pc_when_branch[26]~49 )))) # (!pc_plus_4_M[27] & ((imm_M[15] & (!\pc_when_branch[26]~49 )) # (!imm_M[15] & ((\pc_when_branch[26]~49 ) # 
// (GND)))))
// \pc_when_branch[27]~51  = CARRY((pc_plus_4_M[27] & (!imm_M[15] & !\pc_when_branch[26]~49 )) # (!pc_plus_4_M[27] & ((!\pc_when_branch[26]~49 ) # (!imm_M[15]))))

	.dataa(pc_plus_4_M[27]),
	.datab(imm_M[15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[26]~49 ),
	.combout(\pc_when_branch[27]~50_combout ),
	.cout(\pc_when_branch[27]~51 ));
// synopsys translate_off
defparam \pc_when_branch[27]~50 .lut_mask = 16'h9617;
defparam \pc_when_branch[27]~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X59_Y37_N27
dffeas \rdata1_M[27] (
	.clk(CLK),
	.d(\rdata1_M[27]~25_combout ),
	.asdata(\wdat_WB[27]~11_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[27]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[27] .is_wysiwyg = "true";
defparam \rdata1_M[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N18
cycloneive_lcell_comb \pc_plus_4[26]~48 (
// Equation(s):
// \pc_plus_4[26]~48_combout  = (pc_out_26 & (\pc_plus_4[25]~47  $ (GND))) # (!pc_out_26 & (!\pc_plus_4[25]~47  & VCC))
// \pc_plus_4[26]~49  = CARRY((pc_out_26 & !\pc_plus_4[25]~47 ))

	.dataa(gnd),
	.datab(pc_out_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[25]~47 ),
	.combout(\pc_plus_4[26]~48_combout ),
	.cout(\pc_plus_4[26]~49 ));
// synopsys translate_off
defparam \pc_plus_4[26]~48 .lut_mask = 16'hC30C;
defparam \pc_plus_4[26]~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X59_Y35_N9
dffeas \rdata1_M[26] (
	.clk(CLK),
	.d(\rdata1_M[26]~24_combout ),
	.asdata(\wdat_WB[26]~13_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[26]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[26] .is_wysiwyg = "true";
defparam \rdata1_M[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N22
cycloneive_lcell_comb \pc_plus_4[28]~52 (
// Equation(s):
// \pc_plus_4[28]~52_combout  = (pc_out_28 & (\pc_plus_4[27]~51  $ (GND))) # (!pc_out_28 & (!\pc_plus_4[27]~51  & VCC))
// \pc_plus_4[28]~53  = CARRY((pc_out_28 & !\pc_plus_4[27]~51 ))

	.dataa(pc_out_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[27]~51 ),
	.combout(\pc_plus_4[28]~52_combout ),
	.cout(\pc_plus_4[28]~53 ));
// synopsys translate_off
defparam \pc_plus_4[28]~52 .lut_mask = 16'hA50A;
defparam \pc_plus_4[28]~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N24
cycloneive_lcell_comb \pc_plus_4[29]~54 (
// Equation(s):
// \pc_plus_4[29]~54_combout  = (pc_out_29 & (!\pc_plus_4[28]~53 )) # (!pc_out_29 & ((\pc_plus_4[28]~53 ) # (GND)))
// \pc_plus_4[29]~55  = CARRY((!\pc_plus_4[28]~53 ) # (!pc_out_29))

	.dataa(pc_out_29),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[28]~53 ),
	.combout(\pc_plus_4[29]~54_combout ),
	.cout(\pc_plus_4[29]~55 ));
// synopsys translate_off
defparam \pc_plus_4[29]~54 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[29]~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N22
cycloneive_lcell_comb \pc_when_branch[28]~52 (
// Equation(s):
// \pc_when_branch[28]~52_combout  = ((pc_plus_4_M[28] $ (imm_M[15] $ (!\pc_when_branch[27]~51 )))) # (GND)
// \pc_when_branch[28]~53  = CARRY((pc_plus_4_M[28] & ((imm_M[15]) # (!\pc_when_branch[27]~51 ))) # (!pc_plus_4_M[28] & (imm_M[15] & !\pc_when_branch[27]~51 )))

	.dataa(pc_plus_4_M[28]),
	.datab(imm_M[15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[27]~51 ),
	.combout(\pc_when_branch[28]~52_combout ),
	.cout(\pc_when_branch[28]~53 ));
// synopsys translate_off
defparam \pc_when_branch[28]~52 .lut_mask = 16'h698E;
defparam \pc_when_branch[28]~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N24
cycloneive_lcell_comb \pc_when_branch[29]~54 (
// Equation(s):
// \pc_when_branch[29]~54_combout  = (pc_plus_4_M[29] & ((imm_M[15] & (\pc_when_branch[28]~53  & VCC)) # (!imm_M[15] & (!\pc_when_branch[28]~53 )))) # (!pc_plus_4_M[29] & ((imm_M[15] & (!\pc_when_branch[28]~53 )) # (!imm_M[15] & ((\pc_when_branch[28]~53 ) # 
// (GND)))))
// \pc_when_branch[29]~55  = CARRY((pc_plus_4_M[29] & (!imm_M[15] & !\pc_when_branch[28]~53 )) # (!pc_plus_4_M[29] & ((!\pc_when_branch[28]~53 ) # (!imm_M[15]))))

	.dataa(pc_plus_4_M[29]),
	.datab(imm_M[15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[28]~53 ),
	.combout(\pc_when_branch[29]~54_combout ),
	.cout(\pc_when_branch[29]~55 ));
// synopsys translate_off
defparam \pc_when_branch[29]~54 .lut_mask = 16'h9617;
defparam \pc_when_branch[29]~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X65_Y35_N27
dffeas \rdata1_M[29] (
	.clk(CLK),
	.d(\rdata1_M[29]~27_combout ),
	.asdata(\wdat_WB[29]~7_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[29]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[29] .is_wysiwyg = "true";
defparam \rdata1_M[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y29_N5
dffeas \rdata1_M[28] (
	.clk(CLK),
	.d(\rdata1_M[28]~26_combout ),
	.asdata(\wdat_WB[28]~9_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[28]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[28] .is_wysiwyg = "true";
defparam \rdata1_M[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N26
cycloneive_lcell_comb \pc_plus_4[30]~56 (
// Equation(s):
// \pc_plus_4[30]~56_combout  = (pc_out_30 & (\pc_plus_4[29]~55  $ (GND))) # (!pc_out_30 & (!\pc_plus_4[29]~55  & VCC))
// \pc_plus_4[30]~57  = CARRY((pc_out_30 & !\pc_plus_4[29]~55 ))

	.dataa(pc_out_30),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[29]~55 ),
	.combout(\pc_plus_4[30]~56_combout ),
	.cout(\pc_plus_4[30]~57 ));
// synopsys translate_off
defparam \pc_plus_4[30]~56 .lut_mask = 16'hA50A;
defparam \pc_plus_4[30]~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N28
cycloneive_lcell_comb \pc_plus_4[31]~58 (
// Equation(s):
// \pc_plus_4[31]~58_combout  = \pc_plus_4[30]~57  $ (pc_out_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pc_out_31),
	.cin(\pc_plus_4[30]~57 ),
	.combout(\pc_plus_4[31]~58_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4[31]~58 .lut_mask = 16'h0FF0;
defparam \pc_plus_4[31]~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N26
cycloneive_lcell_comb \pc_when_branch[30]~56 (
// Equation(s):
// \pc_when_branch[30]~56_combout  = ((pc_plus_4_M[30] $ (imm_M[15] $ (!\pc_when_branch[29]~55 )))) # (GND)
// \pc_when_branch[30]~57  = CARRY((pc_plus_4_M[30] & ((imm_M[15]) # (!\pc_when_branch[29]~55 ))) # (!pc_plus_4_M[30] & (imm_M[15] & !\pc_when_branch[29]~55 )))

	.dataa(pc_plus_4_M[30]),
	.datab(imm_M[15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_when_branch[29]~55 ),
	.combout(\pc_when_branch[30]~56_combout ),
	.cout(\pc_when_branch[30]~57 ));
// synopsys translate_off
defparam \pc_when_branch[30]~56 .lut_mask = 16'h698E;
defparam \pc_when_branch[30]~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N28
cycloneive_lcell_comb \pc_when_branch[31]~58 (
// Equation(s):
// \pc_when_branch[31]~58_combout  = pc_plus_4_M[31] $ (\pc_when_branch[30]~57  $ (imm_M[15]))

	.dataa(gnd),
	.datab(pc_plus_4_M[31]),
	.datac(gnd),
	.datad(imm_M[15]),
	.cin(\pc_when_branch[30]~57 ),
	.combout(\pc_when_branch[31]~58_combout ),
	.cout());
// synopsys translate_off
defparam \pc_when_branch[31]~58 .lut_mask = 16'hC33C;
defparam \pc_when_branch[31]~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X65_Y35_N1
dffeas \rdata1_M[31] (
	.clk(CLK),
	.d(\rdata1_M[31]~29_combout ),
	.asdata(\wdat_WB[31]~3_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[31]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[31] .is_wysiwyg = "true";
defparam \rdata1_M[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N15
dffeas \rdata1_M[30] (
	.clk(CLK),
	.d(\rdata1_M[30]~28_combout ),
	.asdata(\wdat_WB[30]~5_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(\rdata1_M~33_combout ),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_M[30]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_M[30] .is_wysiwyg = "true";
defparam \rdata1_M[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N2
cycloneive_lcell_comb \Add2~0 (
// Equation(s):
// \Add2~0_combout  = pc_plus_4_M[2] $ (VCC)
// \Add2~1  = CARRY(pc_plus_4_M[2])

	.dataa(gnd),
	.datab(pc_plus_4_M[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout(\Add2~1 ));
// synopsys translate_off
defparam \Add2~0 .lut_mask = 16'h33CC;
defparam \Add2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N4
cycloneive_lcell_comb \Add2~2 (
// Equation(s):
// \Add2~2_combout  = (pc_plus_4_M[3] & (\Add2~1  & VCC)) # (!pc_plus_4_M[3] & (!\Add2~1 ))
// \Add2~3  = CARRY((!pc_plus_4_M[3] & !\Add2~1 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~1 ),
	.combout(\Add2~2_combout ),
	.cout(\Add2~3 ));
// synopsys translate_off
defparam \Add2~2 .lut_mask = 16'hC303;
defparam \Add2~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N6
cycloneive_lcell_comb \Add2~4 (
// Equation(s):
// \Add2~4_combout  = (pc_plus_4_M[4] & ((GND) # (!\Add2~3 ))) # (!pc_plus_4_M[4] & (\Add2~3  $ (GND)))
// \Add2~5  = CARRY((pc_plus_4_M[4]) # (!\Add2~3 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~3 ),
	.combout(\Add2~4_combout ),
	.cout(\Add2~5 ));
// synopsys translate_off
defparam \Add2~4 .lut_mask = 16'h3CCF;
defparam \Add2~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N8
cycloneive_lcell_comb \Add2~6 (
// Equation(s):
// \Add2~6_combout  = (pc_plus_4_M[5] & (\Add2~5  & VCC)) # (!pc_plus_4_M[5] & (!\Add2~5 ))
// \Add2~7  = CARRY((!pc_plus_4_M[5] & !\Add2~5 ))

	.dataa(pc_plus_4_M[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~5 ),
	.combout(\Add2~6_combout ),
	.cout(\Add2~7 ));
// synopsys translate_off
defparam \Add2~6 .lut_mask = 16'hA505;
defparam \Add2~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N10
cycloneive_lcell_comb \Add2~8 (
// Equation(s):
// \Add2~8_combout  = (pc_plus_4_M[6] & ((GND) # (!\Add2~7 ))) # (!pc_plus_4_M[6] & (\Add2~7  $ (GND)))
// \Add2~9  = CARRY((pc_plus_4_M[6]) # (!\Add2~7 ))

	.dataa(pc_plus_4_M[6]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~7 ),
	.combout(\Add2~8_combout ),
	.cout(\Add2~9 ));
// synopsys translate_off
defparam \Add2~8 .lut_mask = 16'h5AAF;
defparam \Add2~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N12
cycloneive_lcell_comb \Add2~10 (
// Equation(s):
// \Add2~10_combout  = (pc_plus_4_M[7] & (\Add2~9  & VCC)) # (!pc_plus_4_M[7] & (!\Add2~9 ))
// \Add2~11  = CARRY((!pc_plus_4_M[7] & !\Add2~9 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[7]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~9 ),
	.combout(\Add2~10_combout ),
	.cout(\Add2~11 ));
// synopsys translate_off
defparam \Add2~10 .lut_mask = 16'hC303;
defparam \Add2~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N14
cycloneive_lcell_comb \Add2~12 (
// Equation(s):
// \Add2~12_combout  = (pc_plus_4_M[8] & ((GND) # (!\Add2~11 ))) # (!pc_plus_4_M[8] & (\Add2~11  $ (GND)))
// \Add2~13  = CARRY((pc_plus_4_M[8]) # (!\Add2~11 ))

	.dataa(pc_plus_4_M[8]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~11 ),
	.combout(\Add2~12_combout ),
	.cout(\Add2~13 ));
// synopsys translate_off
defparam \Add2~12 .lut_mask = 16'h5AAF;
defparam \Add2~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N16
cycloneive_lcell_comb \Add2~14 (
// Equation(s):
// \Add2~14_combout  = (pc_plus_4_M[9] & (\Add2~13  & VCC)) # (!pc_plus_4_M[9] & (!\Add2~13 ))
// \Add2~15  = CARRY((!pc_plus_4_M[9] & !\Add2~13 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[9]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~13 ),
	.combout(\Add2~14_combout ),
	.cout(\Add2~15 ));
// synopsys translate_off
defparam \Add2~14 .lut_mask = 16'hC303;
defparam \Add2~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N18
cycloneive_lcell_comb \Add2~16 (
// Equation(s):
// \Add2~16_combout  = (pc_plus_4_M[10] & ((GND) # (!\Add2~15 ))) # (!pc_plus_4_M[10] & (\Add2~15  $ (GND)))
// \Add2~17  = CARRY((pc_plus_4_M[10]) # (!\Add2~15 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[10]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~15 ),
	.combout(\Add2~16_combout ),
	.cout(\Add2~17 ));
// synopsys translate_off
defparam \Add2~16 .lut_mask = 16'h3CCF;
defparam \Add2~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N20
cycloneive_lcell_comb \Add2~18 (
// Equation(s):
// \Add2~18_combout  = (pc_plus_4_M[11] & (\Add2~17  & VCC)) # (!pc_plus_4_M[11] & (!\Add2~17 ))
// \Add2~19  = CARRY((!pc_plus_4_M[11] & !\Add2~17 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[11]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~17 ),
	.combout(\Add2~18_combout ),
	.cout(\Add2~19 ));
// synopsys translate_off
defparam \Add2~18 .lut_mask = 16'hC303;
defparam \Add2~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N22
cycloneive_lcell_comb \Add2~20 (
// Equation(s):
// \Add2~20_combout  = (pc_plus_4_M[12] & ((GND) # (!\Add2~19 ))) # (!pc_plus_4_M[12] & (\Add2~19  $ (GND)))
// \Add2~21  = CARRY((pc_plus_4_M[12]) # (!\Add2~19 ))

	.dataa(pc_plus_4_M[12]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~19 ),
	.combout(\Add2~20_combout ),
	.cout(\Add2~21 ));
// synopsys translate_off
defparam \Add2~20 .lut_mask = 16'h5AAF;
defparam \Add2~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N24
cycloneive_lcell_comb \Add2~22 (
// Equation(s):
// \Add2~22_combout  = (pc_plus_4_M[13] & (\Add2~21  & VCC)) # (!pc_plus_4_M[13] & (!\Add2~21 ))
// \Add2~23  = CARRY((!pc_plus_4_M[13] & !\Add2~21 ))

	.dataa(pc_plus_4_M[13]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~21 ),
	.combout(\Add2~22_combout ),
	.cout(\Add2~23 ));
// synopsys translate_off
defparam \Add2~22 .lut_mask = 16'hA505;
defparam \Add2~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N26
cycloneive_lcell_comb \Add2~24 (
// Equation(s):
// \Add2~24_combout  = (pc_plus_4_M[14] & ((GND) # (!\Add2~23 ))) # (!pc_plus_4_M[14] & (\Add2~23  $ (GND)))
// \Add2~25  = CARRY((pc_plus_4_M[14]) # (!\Add2~23 ))

	.dataa(pc_plus_4_M[14]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~23 ),
	.combout(\Add2~24_combout ),
	.cout(\Add2~25 ));
// synopsys translate_off
defparam \Add2~24 .lut_mask = 16'h5AAF;
defparam \Add2~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N28
cycloneive_lcell_comb \Add2~26 (
// Equation(s):
// \Add2~26_combout  = (pc_plus_4_M[15] & (\Add2~25  & VCC)) # (!pc_plus_4_M[15] & (!\Add2~25 ))
// \Add2~27  = CARRY((!pc_plus_4_M[15] & !\Add2~25 ))

	.dataa(pc_plus_4_M[15]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~25 ),
	.combout(\Add2~26_combout ),
	.cout(\Add2~27 ));
// synopsys translate_off
defparam \Add2~26 .lut_mask = 16'hA505;
defparam \Add2~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N30
cycloneive_lcell_comb \Add2~28 (
// Equation(s):
// \Add2~28_combout  = (pc_plus_4_M[16] & ((GND) # (!\Add2~27 ))) # (!pc_plus_4_M[16] & (\Add2~27  $ (GND)))
// \Add2~29  = CARRY((pc_plus_4_M[16]) # (!\Add2~27 ))

	.dataa(pc_plus_4_M[16]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~27 ),
	.combout(\Add2~28_combout ),
	.cout(\Add2~29 ));
// synopsys translate_off
defparam \Add2~28 .lut_mask = 16'h5AAF;
defparam \Add2~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N0
cycloneive_lcell_comb \Add2~30 (
// Equation(s):
// \Add2~30_combout  = (pc_plus_4_M[17] & (\Add2~29  & VCC)) # (!pc_plus_4_M[17] & (!\Add2~29 ))
// \Add2~31  = CARRY((!pc_plus_4_M[17] & !\Add2~29 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[17]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~29 ),
	.combout(\Add2~30_combout ),
	.cout(\Add2~31 ));
// synopsys translate_off
defparam \Add2~30 .lut_mask = 16'hC303;
defparam \Add2~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N2
cycloneive_lcell_comb \Add2~32 (
// Equation(s):
// \Add2~32_combout  = (pc_plus_4_M[18] & ((GND) # (!\Add2~31 ))) # (!pc_plus_4_M[18] & (\Add2~31  $ (GND)))
// \Add2~33  = CARRY((pc_plus_4_M[18]) # (!\Add2~31 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[18]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~31 ),
	.combout(\Add2~32_combout ),
	.cout(\Add2~33 ));
// synopsys translate_off
defparam \Add2~32 .lut_mask = 16'h3CCF;
defparam \Add2~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N4
cycloneive_lcell_comb \Add2~34 (
// Equation(s):
// \Add2~34_combout  = (pc_plus_4_M[19] & (\Add2~33  & VCC)) # (!pc_plus_4_M[19] & (!\Add2~33 ))
// \Add2~35  = CARRY((!pc_plus_4_M[19] & !\Add2~33 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[19]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~33 ),
	.combout(\Add2~34_combout ),
	.cout(\Add2~35 ));
// synopsys translate_off
defparam \Add2~34 .lut_mask = 16'hC303;
defparam \Add2~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N6
cycloneive_lcell_comb \Add2~36 (
// Equation(s):
// \Add2~36_combout  = (pc_plus_4_M[20] & ((GND) # (!\Add2~35 ))) # (!pc_plus_4_M[20] & (\Add2~35  $ (GND)))
// \Add2~37  = CARRY((pc_plus_4_M[20]) # (!\Add2~35 ))

	.dataa(pc_plus_4_M[20]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~35 ),
	.combout(\Add2~36_combout ),
	.cout(\Add2~37 ));
// synopsys translate_off
defparam \Add2~36 .lut_mask = 16'h5AAF;
defparam \Add2~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N8
cycloneive_lcell_comb \Add2~38 (
// Equation(s):
// \Add2~38_combout  = (pc_plus_4_M[21] & (\Add2~37  & VCC)) # (!pc_plus_4_M[21] & (!\Add2~37 ))
// \Add2~39  = CARRY((!pc_plus_4_M[21] & !\Add2~37 ))

	.dataa(pc_plus_4_M[21]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~37 ),
	.combout(\Add2~38_combout ),
	.cout(\Add2~39 ));
// synopsys translate_off
defparam \Add2~38 .lut_mask = 16'hA505;
defparam \Add2~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N10
cycloneive_lcell_comb \Add2~40 (
// Equation(s):
// \Add2~40_combout  = (pc_plus_4_M[22] & ((GND) # (!\Add2~39 ))) # (!pc_plus_4_M[22] & (\Add2~39  $ (GND)))
// \Add2~41  = CARRY((pc_plus_4_M[22]) # (!\Add2~39 ))

	.dataa(pc_plus_4_M[22]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~39 ),
	.combout(\Add2~40_combout ),
	.cout(\Add2~41 ));
// synopsys translate_off
defparam \Add2~40 .lut_mask = 16'h5AAF;
defparam \Add2~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N12
cycloneive_lcell_comb \Add2~42 (
// Equation(s):
// \Add2~42_combout  = (pc_plus_4_M[23] & (\Add2~41  & VCC)) # (!pc_plus_4_M[23] & (!\Add2~41 ))
// \Add2~43  = CARRY((!pc_plus_4_M[23] & !\Add2~41 ))

	.dataa(pc_plus_4_M[23]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~41 ),
	.combout(\Add2~42_combout ),
	.cout(\Add2~43 ));
// synopsys translate_off
defparam \Add2~42 .lut_mask = 16'hA505;
defparam \Add2~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N14
cycloneive_lcell_comb \Add2~44 (
// Equation(s):
// \Add2~44_combout  = (pc_plus_4_M[24] & ((GND) # (!\Add2~43 ))) # (!pc_plus_4_M[24] & (\Add2~43  $ (GND)))
// \Add2~45  = CARRY((pc_plus_4_M[24]) # (!\Add2~43 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[24]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~43 ),
	.combout(\Add2~44_combout ),
	.cout(\Add2~45 ));
// synopsys translate_off
defparam \Add2~44 .lut_mask = 16'h3CCF;
defparam \Add2~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N16
cycloneive_lcell_comb \Add2~46 (
// Equation(s):
// \Add2~46_combout  = (pc_plus_4_M[25] & (\Add2~45  & VCC)) # (!pc_plus_4_M[25] & (!\Add2~45 ))
// \Add2~47  = CARRY((!pc_plus_4_M[25] & !\Add2~45 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[25]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~45 ),
	.combout(\Add2~46_combout ),
	.cout(\Add2~47 ));
// synopsys translate_off
defparam \Add2~46 .lut_mask = 16'hC303;
defparam \Add2~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N18
cycloneive_lcell_comb \Add2~48 (
// Equation(s):
// \Add2~48_combout  = (pc_plus_4_M[26] & ((GND) # (!\Add2~47 ))) # (!pc_plus_4_M[26] & (\Add2~47  $ (GND)))
// \Add2~49  = CARRY((pc_plus_4_M[26]) # (!\Add2~47 ))

	.dataa(pc_plus_4_M[26]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~47 ),
	.combout(\Add2~48_combout ),
	.cout(\Add2~49 ));
// synopsys translate_off
defparam \Add2~48 .lut_mask = 16'h5AAF;
defparam \Add2~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N20
cycloneive_lcell_comb \Add2~50 (
// Equation(s):
// \Add2~50_combout  = (pc_plus_4_M[27] & (\Add2~49  & VCC)) # (!pc_plus_4_M[27] & (!\Add2~49 ))
// \Add2~51  = CARRY((!pc_plus_4_M[27] & !\Add2~49 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[27]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~49 ),
	.combout(\Add2~50_combout ),
	.cout(\Add2~51 ));
// synopsys translate_off
defparam \Add2~50 .lut_mask = 16'hC303;
defparam \Add2~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N22
cycloneive_lcell_comb \Add2~52 (
// Equation(s):
// \Add2~52_combout  = (pc_plus_4_M[28] & ((GND) # (!\Add2~51 ))) # (!pc_plus_4_M[28] & (\Add2~51  $ (GND)))
// \Add2~53  = CARRY((pc_plus_4_M[28]) # (!\Add2~51 ))

	.dataa(pc_plus_4_M[28]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~51 ),
	.combout(\Add2~52_combout ),
	.cout(\Add2~53 ));
// synopsys translate_off
defparam \Add2~52 .lut_mask = 16'h5AAF;
defparam \Add2~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N24
cycloneive_lcell_comb \Add2~54 (
// Equation(s):
// \Add2~54_combout  = (pc_plus_4_M[29] & (\Add2~53  & VCC)) # (!pc_plus_4_M[29] & (!\Add2~53 ))
// \Add2~55  = CARRY((!pc_plus_4_M[29] & !\Add2~53 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[29]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~53 ),
	.combout(\Add2~54_combout ),
	.cout(\Add2~55 ));
// synopsys translate_off
defparam \Add2~54 .lut_mask = 16'hC303;
defparam \Add2~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N26
cycloneive_lcell_comb \Add2~56 (
// Equation(s):
// \Add2~56_combout  = (pc_plus_4_M[30] & ((GND) # (!\Add2~55 ))) # (!pc_plus_4_M[30] & (\Add2~55  $ (GND)))
// \Add2~57  = CARRY((pc_plus_4_M[30]) # (!\Add2~55 ))

	.dataa(gnd),
	.datab(pc_plus_4_M[30]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~55 ),
	.combout(\Add2~56_combout ),
	.cout(\Add2~57 ));
// synopsys translate_off
defparam \Add2~56 .lut_mask = 16'h3CCF;
defparam \Add2~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N28
cycloneive_lcell_comb \Add2~58 (
// Equation(s):
// \Add2~58_combout  = \Add2~57  $ (!pc_plus_4_M[31])

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pc_plus_4_M[31]),
	.cin(\Add2~57 ),
	.combout(\Add2~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add2~58 .lut_mask = 16'hF00F;
defparam \Add2~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N12
cycloneive_lcell_comb \rdata1_M[1]~31 (
// Equation(s):
// \rdata1_M[1]~31_combout  = (\rdata1_M~32_combout  & ((porto_M_1))) # (!\rdata1_M~32_combout  & (rdata1_EX[1]))

	.dataa(rdata1_EX[1]),
	.datab(porto_M_1),
	.datac(gnd),
	.datad(\rdata1_M~32_combout ),
	.cin(gnd),
	.combout(\rdata1_M[1]~31_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[1]~31 .lut_mask = 16'hCCAA;
defparam \rdata1_M[1]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N22
cycloneive_lcell_comb \rdata1_M[0]~30 (
// Equation(s):
// \rdata1_M[0]~30_combout  = (\rdata1_M~32_combout  & (porto_M_0)) # (!\rdata1_M~32_combout  & ((rdata1_EX[0])))

	.dataa(porto_M_0),
	.datab(rdata1_EX[0]),
	.datac(gnd),
	.datad(\rdata1_M~32_combout ),
	.cin(gnd),
	.combout(\rdata1_M[0]~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[0]~30 .lut_mask = 16'hAACC;
defparam \rdata1_M[0]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N28
cycloneive_lcell_comb \rdata1_M[3]~0 (
// Equation(s):
// \rdata1_M[3]~0_combout  = (\rdata1_M~32_combout  & ((porto_M_3))) # (!\rdata1_M~32_combout  & (rdata1_EX[3]))

	.dataa(\rdata1_M~32_combout ),
	.datab(rdata1_EX[3]),
	.datac(gnd),
	.datad(porto_M_3),
	.cin(gnd),
	.combout(\rdata1_M[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[3]~0 .lut_mask = 16'hEE44;
defparam \rdata1_M[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N24
cycloneive_lcell_comb \rdata1_M[2]~1 (
// Equation(s):
// \rdata1_M[2]~1_combout  = (\rdata1_M~32_combout  & (porto_M_2)) # (!\rdata1_M~32_combout  & ((rdata1_EX[2])))

	.dataa(porto_M_2),
	.datab(\rdata1_M~32_combout ),
	.datac(gnd),
	.datad(rdata1_EX[2]),
	.cin(gnd),
	.combout(\rdata1_M[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[2]~1 .lut_mask = 16'hBB88;
defparam \rdata1_M[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N28
cycloneive_lcell_comb \rdata1_M[5]~3 (
// Equation(s):
// \rdata1_M[5]~3_combout  = (\rdata1_M~32_combout  & ((porto_M_5))) # (!\rdata1_M~32_combout  & (rdata1_EX[5]))

	.dataa(\rdata1_M~32_combout ),
	.datab(rdata1_EX[5]),
	.datac(gnd),
	.datad(porto_M_5),
	.cin(gnd),
	.combout(\rdata1_M[5]~3_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[5]~3 .lut_mask = 16'hEE44;
defparam \rdata1_M[5]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N6
cycloneive_lcell_comb \rdata1_M[4]~2 (
// Equation(s):
// \rdata1_M[4]~2_combout  = (\rdata1_M~32_combout  & (porto_M_4)) # (!\rdata1_M~32_combout  & ((rdata1_EX[4])))

	.dataa(\rdata1_M~32_combout ),
	.datab(porto_M_4),
	.datac(gnd),
	.datad(rdata1_EX[4]),
	.cin(gnd),
	.combout(\rdata1_M[4]~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[4]~2 .lut_mask = 16'hDD88;
defparam \rdata1_M[4]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N12
cycloneive_lcell_comb \rdata1_M[7]~5 (
// Equation(s):
// \rdata1_M[7]~5_combout  = (\rdata1_M~32_combout  & ((porto_M_7))) # (!\rdata1_M~32_combout  & (rdata1_EX[7]))

	.dataa(\rdata1_M~32_combout ),
	.datab(rdata1_EX[7]),
	.datac(gnd),
	.datad(porto_M_7),
	.cin(gnd),
	.combout(\rdata1_M[7]~5_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[7]~5 .lut_mask = 16'hEE44;
defparam \rdata1_M[7]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N8
cycloneive_lcell_comb \rdata1_M[6]~4 (
// Equation(s):
// \rdata1_M[6]~4_combout  = (\rdata1_M~32_combout  & ((porto_M_6))) # (!\rdata1_M~32_combout  & (rdata1_EX[6]))

	.dataa(rdata1_EX[6]),
	.datab(porto_M_6),
	.datac(gnd),
	.datad(\rdata1_M~32_combout ),
	.cin(gnd),
	.combout(\rdata1_M[6]~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[6]~4 .lut_mask = 16'hCCAA;
defparam \rdata1_M[6]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N2
cycloneive_lcell_comb \rdata1_M[9]~7 (
// Equation(s):
// \rdata1_M[9]~7_combout  = (\rdata1_M~32_combout  & (porto_M_9)) # (!\rdata1_M~32_combout  & ((rdata1_EX[9])))

	.dataa(\rdata1_M~32_combout ),
	.datab(porto_M_9),
	.datac(gnd),
	.datad(rdata1_EX[9]),
	.cin(gnd),
	.combout(\rdata1_M[9]~7_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[9]~7 .lut_mask = 16'hDD88;
defparam \rdata1_M[9]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N24
cycloneive_lcell_comb \rdata1_M[8]~6 (
// Equation(s):
// \rdata1_M[8]~6_combout  = (\rdata1_M~32_combout  & ((porto_M_8))) # (!\rdata1_M~32_combout  & (rdata1_EX[8]))

	.dataa(rdata1_EX[8]),
	.datab(porto_M_8),
	.datac(gnd),
	.datad(\rdata1_M~32_combout ),
	.cin(gnd),
	.combout(\rdata1_M[8]~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[8]~6 .lut_mask = 16'hCCAA;
defparam \rdata1_M[8]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N0
cycloneive_lcell_comb \rdata1_M[11]~9 (
// Equation(s):
// \rdata1_M[11]~9_combout  = (\rdata1_M~32_combout  & ((porto_M_11))) # (!\rdata1_M~32_combout  & (rdata1_EX[11]))

	.dataa(\rdata1_M~32_combout ),
	.datab(rdata1_EX[11]),
	.datac(gnd),
	.datad(porto_M_11),
	.cin(gnd),
	.combout(\rdata1_M[11]~9_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[11]~9 .lut_mask = 16'hEE44;
defparam \rdata1_M[11]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N12
cycloneive_lcell_comb \rdata1_M[10]~8 (
// Equation(s):
// \rdata1_M[10]~8_combout  = (\rdata1_M~32_combout  & (porto_M_10)) # (!\rdata1_M~32_combout  & ((rdata1_EX[10])))

	.dataa(porto_M_10),
	.datab(rdata1_EX[10]),
	.datac(gnd),
	.datad(\rdata1_M~32_combout ),
	.cin(gnd),
	.combout(\rdata1_M[10]~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[10]~8 .lut_mask = 16'hAACC;
defparam \rdata1_M[10]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N4
cycloneive_lcell_comb \rdata1_M[13]~11 (
// Equation(s):
// \rdata1_M[13]~11_combout  = (\rdata1_M~32_combout  & ((porto_M_13))) # (!\rdata1_M~32_combout  & (rdata1_EX[13]))

	.dataa(\rdata1_M~32_combout ),
	.datab(rdata1_EX[13]),
	.datac(gnd),
	.datad(porto_M_13),
	.cin(gnd),
	.combout(\rdata1_M[13]~11_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[13]~11 .lut_mask = 16'hEE44;
defparam \rdata1_M[13]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N28
cycloneive_lcell_comb \rdata1_M[12]~10 (
// Equation(s):
// \rdata1_M[12]~10_combout  = (\rdata1_M~32_combout  & ((porto_M_12))) # (!\rdata1_M~32_combout  & (rdata1_EX[12]))

	.dataa(rdata1_EX[12]),
	.datab(porto_M_12),
	.datac(gnd),
	.datad(\rdata1_M~32_combout ),
	.cin(gnd),
	.combout(\rdata1_M[12]~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[12]~10 .lut_mask = 16'hCCAA;
defparam \rdata1_M[12]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N26
cycloneive_lcell_comb \rdata1_M[15]~13 (
// Equation(s):
// \rdata1_M[15]~13_combout  = (\rdata1_M~32_combout  & (porto_M_15)) # (!\rdata1_M~32_combout  & ((rdata1_EX[15])))

	.dataa(\rdata1_M~32_combout ),
	.datab(porto_M_15),
	.datac(gnd),
	.datad(rdata1_EX[15]),
	.cin(gnd),
	.combout(\rdata1_M[15]~13_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[15]~13 .lut_mask = 16'hDD88;
defparam \rdata1_M[15]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N16
cycloneive_lcell_comb \rdata1_M[14]~12 (
// Equation(s):
// \rdata1_M[14]~12_combout  = (\rdata1_M~32_combout  & ((porto_M_14))) # (!\rdata1_M~32_combout  & (rdata1_EX[14]))

	.dataa(\rdata1_M~32_combout ),
	.datab(rdata1_EX[14]),
	.datac(gnd),
	.datad(porto_M_14),
	.cin(gnd),
	.combout(\rdata1_M[14]~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[14]~12 .lut_mask = 16'hEE44;
defparam \rdata1_M[14]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N2
cycloneive_lcell_comb \rdata1_M[17]~15 (
// Equation(s):
// \rdata1_M[17]~15_combout  = (\rdata1_M~32_combout  & ((porto_M_17))) # (!\rdata1_M~32_combout  & (rdata1_EX[17]))

	.dataa(\rdata1_M~32_combout ),
	.datab(rdata1_EX[17]),
	.datac(gnd),
	.datad(porto_M_17),
	.cin(gnd),
	.combout(\rdata1_M[17]~15_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[17]~15 .lut_mask = 16'hEE44;
defparam \rdata1_M[17]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N22
cycloneive_lcell_comb \rdata1_M[16]~14 (
// Equation(s):
// \rdata1_M[16]~14_combout  = (\rdata1_M~32_combout  & (porto_M_16)) # (!\rdata1_M~32_combout  & ((rdata1_EX[16])))

	.dataa(porto_M_16),
	.datab(rdata1_EX[16]),
	.datac(gnd),
	.datad(\rdata1_M~32_combout ),
	.cin(gnd),
	.combout(\rdata1_M[16]~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[16]~14 .lut_mask = 16'hAACC;
defparam \rdata1_M[16]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N10
cycloneive_lcell_comb \rdata1_M[19]~17 (
// Equation(s):
// \rdata1_M[19]~17_combout  = (\rdata1_M~32_combout  & ((porto_M_19))) # (!\rdata1_M~32_combout  & (rdata1_EX[19]))

	.dataa(rdata1_EX[19]),
	.datab(\rdata1_M~32_combout ),
	.datac(gnd),
	.datad(porto_M_19),
	.cin(gnd),
	.combout(\rdata1_M[19]~17_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[19]~17 .lut_mask = 16'hEE22;
defparam \rdata1_M[19]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N0
cycloneive_lcell_comb \rdata1_M[18]~16 (
// Equation(s):
// \rdata1_M[18]~16_combout  = (\rdata1_M~32_combout  & ((porto_M_18))) # (!\rdata1_M~32_combout  & (rdata1_EX[18]))

	.dataa(\rdata1_M~32_combout ),
	.datab(rdata1_EX[18]),
	.datac(gnd),
	.datad(porto_M_18),
	.cin(gnd),
	.combout(\rdata1_M[18]~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[18]~16 .lut_mask = 16'hEE44;
defparam \rdata1_M[18]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N26
cycloneive_lcell_comb \rdata1_M[21]~19 (
// Equation(s):
// \rdata1_M[21]~19_combout  = (\rdata1_M~32_combout  & (porto_M_21)) # (!\rdata1_M~32_combout  & ((rdata1_EX[21])))

	.dataa(porto_M_21),
	.datab(\rdata1_M~32_combout ),
	.datac(gnd),
	.datad(rdata1_EX[21]),
	.cin(gnd),
	.combout(\rdata1_M[21]~19_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[21]~19 .lut_mask = 16'hBB88;
defparam \rdata1_M[21]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N8
cycloneive_lcell_comb \rdata1_M[20]~18 (
// Equation(s):
// \rdata1_M[20]~18_combout  = (\rdata1_M~32_combout  & (porto_M_20)) # (!\rdata1_M~32_combout  & ((rdata1_EX[20])))

	.dataa(porto_M_20),
	.datab(rdata1_EX[20]),
	.datac(gnd),
	.datad(\rdata1_M~32_combout ),
	.cin(gnd),
	.combout(\rdata1_M[20]~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[20]~18 .lut_mask = 16'hAACC;
defparam \rdata1_M[20]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N24
cycloneive_lcell_comb \rdata1_M[23]~21 (
// Equation(s):
// \rdata1_M[23]~21_combout  = (\rdata1_M~32_combout  & ((porto_M_23))) # (!\rdata1_M~32_combout  & (rdata1_EX[23]))

	.dataa(\rdata1_M~32_combout ),
	.datab(rdata1_EX[23]),
	.datac(gnd),
	.datad(porto_M_23),
	.cin(gnd),
	.combout(\rdata1_M[23]~21_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[23]~21 .lut_mask = 16'hEE44;
defparam \rdata1_M[23]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N10
cycloneive_lcell_comb \rdata1_M[22]~20 (
// Equation(s):
// \rdata1_M[22]~20_combout  = (\rdata1_M~32_combout  & (porto_M_22)) # (!\rdata1_M~32_combout  & ((rdata1_EX[22])))

	.dataa(porto_M_22),
	.datab(\rdata1_M~32_combout ),
	.datac(gnd),
	.datad(rdata1_EX[22]),
	.cin(gnd),
	.combout(\rdata1_M[22]~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[22]~20 .lut_mask = 16'hBB88;
defparam \rdata1_M[22]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N0
cycloneive_lcell_comb \rdata1_M[25]~23 (
// Equation(s):
// \rdata1_M[25]~23_combout  = (\rdata1_M~32_combout  & ((porto_M_25))) # (!\rdata1_M~32_combout  & (rdata1_EX[25]))

	.dataa(rdata1_EX[25]),
	.datab(porto_M_25),
	.datac(gnd),
	.datad(\rdata1_M~32_combout ),
	.cin(gnd),
	.combout(\rdata1_M[25]~23_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[25]~23 .lut_mask = 16'hCCAA;
defparam \rdata1_M[25]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N12
cycloneive_lcell_comb \rdata1_M[24]~22 (
// Equation(s):
// \rdata1_M[24]~22_combout  = (\rdata1_M~32_combout  & ((porto_M_24))) # (!\rdata1_M~32_combout  & (rdata1_EX[24]))

	.dataa(rdata1_EX[24]),
	.datab(porto_M_24),
	.datac(gnd),
	.datad(\rdata1_M~32_combout ),
	.cin(gnd),
	.combout(\rdata1_M[24]~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[24]~22 .lut_mask = 16'hCCAA;
defparam \rdata1_M[24]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N26
cycloneive_lcell_comb \rdata1_M[27]~25 (
// Equation(s):
// \rdata1_M[27]~25_combout  = (\rdata1_M~32_combout  & (porto_M_27)) # (!\rdata1_M~32_combout  & ((rdata1_EX[27])))

	.dataa(porto_M_27),
	.datab(\rdata1_M~32_combout ),
	.datac(gnd),
	.datad(rdata1_EX[27]),
	.cin(gnd),
	.combout(\rdata1_M[27]~25_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[27]~25 .lut_mask = 16'hBB88;
defparam \rdata1_M[27]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N8
cycloneive_lcell_comb \rdata1_M[26]~24 (
// Equation(s):
// \rdata1_M[26]~24_combout  = (\rdata1_M~32_combout  & (porto_M_26)) # (!\rdata1_M~32_combout  & ((rdata1_EX[26])))

	.dataa(porto_M_26),
	.datab(\rdata1_M~32_combout ),
	.datac(gnd),
	.datad(rdata1_EX[26]),
	.cin(gnd),
	.combout(\rdata1_M[26]~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[26]~24 .lut_mask = 16'hBB88;
defparam \rdata1_M[26]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N26
cycloneive_lcell_comb \rdata1_M[29]~27 (
// Equation(s):
// \rdata1_M[29]~27_combout  = (\rdata1_M~32_combout  & ((porto_M_29))) # (!\rdata1_M~32_combout  & (rdata1_EX[29]))

	.dataa(rdata1_EX[29]),
	.datab(\rdata1_M~32_combout ),
	.datac(gnd),
	.datad(porto_M_29),
	.cin(gnd),
	.combout(\rdata1_M[29]~27_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[29]~27 .lut_mask = 16'hEE22;
defparam \rdata1_M[29]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N4
cycloneive_lcell_comb \rdata1_M[28]~26 (
// Equation(s):
// \rdata1_M[28]~26_combout  = (\rdata1_M~32_combout  & (porto_M_28)) # (!\rdata1_M~32_combout  & ((rdata1_EX[28])))

	.dataa(porto_M_28),
	.datab(\rdata1_M~32_combout ),
	.datac(gnd),
	.datad(rdata1_EX[28]),
	.cin(gnd),
	.combout(\rdata1_M[28]~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[28]~26 .lut_mask = 16'hBB88;
defparam \rdata1_M[28]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N0
cycloneive_lcell_comb \rdata1_M[31]~29 (
// Equation(s):
// \rdata1_M[31]~29_combout  = (\rdata1_M~32_combout  & ((porto_M_31))) # (!\rdata1_M~32_combout  & (rdata1_EX[31]))

	.dataa(rdata1_EX[31]),
	.datab(\rdata1_M~32_combout ),
	.datac(gnd),
	.datad(porto_M_31),
	.cin(gnd),
	.combout(\rdata1_M[31]~29_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[31]~29 .lut_mask = 16'hEE22;
defparam \rdata1_M[31]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N14
cycloneive_lcell_comb \rdata1_M[30]~28 (
// Equation(s):
// \rdata1_M[30]~28_combout  = (\rdata1_M~32_combout  & (porto_M_30)) # (!\rdata1_M~32_combout  & ((rdata1_EX[30])))

	.dataa(porto_M_30),
	.datab(\rdata1_M~32_combout ),
	.datac(gnd),
	.datad(rdata1_EX[30]),
	.cin(gnd),
	.combout(\rdata1_M[30]~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M[30]~28 .lut_mask = 16'hBB88;
defparam \rdata1_M[30]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N1
dffeas bne_M(
	.clk(CLK),
	.d(\bne_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bne_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam bne_M.is_wysiwyg = "true";
defparam bne_M.power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N7
dffeas jr_M(
	.clk(CLK),
	.d(\jr_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\jr_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam jr_M.is_wysiwyg = "true";
defparam jr_M.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N5
dffeas \op_EX[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\op_EX~0_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_EX[5]),
	.prn(vcc));
// synopsys translate_off
defparam \op_EX[5] .is_wysiwyg = "true";
defparam \op_EX[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N11
dffeas \op_EX[4] (
	.clk(CLK),
	.d(\op_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_EX[4]),
	.prn(vcc));
// synopsys translate_off
defparam \op_EX[4] .is_wysiwyg = "true";
defparam \op_EX[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N17
dffeas \op_EX[3] (
	.clk(CLK),
	.d(\op_EX~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_EX[3]),
	.prn(vcc));
// synopsys translate_off
defparam \op_EX[3] .is_wysiwyg = "true";
defparam \op_EX[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N7
dffeas \op_EX[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\op_EX~3_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_EX[2]),
	.prn(vcc));
// synopsys translate_off
defparam \op_EX[2] .is_wysiwyg = "true";
defparam \op_EX[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N6
cycloneive_lcell_comb \Equal4~0 (
// Equation(s):
// \Equal4~0_combout  = (op_EX[4] & (op_EX[5] & (op_EX[2] & op_EX[3])))

	.dataa(op_EX[4]),
	.datab(op_EX[5]),
	.datac(op_EX[2]),
	.datad(op_EX[3]),
	.cin(gnd),
	.combout(\Equal4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~0 .lut_mask = 16'h8000;
defparam \Equal4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N23
dffeas \op_EX[1] (
	.clk(CLK),
	.d(\op_EX~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_EX[1]),
	.prn(vcc));
// synopsys translate_off
defparam \op_EX[1] .is_wysiwyg = "true";
defparam \op_EX[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N1
dffeas \op_EX[0] (
	.clk(CLK),
	.d(\op_EX~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_EX[0]),
	.prn(vcc));
// synopsys translate_off
defparam \op_EX[0] .is_wysiwyg = "true";
defparam \op_EX[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N30
cycloneive_lcell_comb \Equal4~1 (
// Equation(s):
// \Equal4~1_combout  = (op_EX[1] & op_EX[0])

	.dataa(gnd),
	.datab(gnd),
	.datac(op_EX[1]),
	.datad(op_EX[0]),
	.cin(gnd),
	.combout(\Equal4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~1 .lut_mask = 16'hF000;
defparam \Equal4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N17
dffeas \instruction_EX[16] (
	.clk(CLK),
	.d(\instruction_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_EX[16]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_EX[16] .is_wysiwyg = "true";
defparam \instruction_EX[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N31
dffeas \instruction_EX[17] (
	.clk(CLK),
	.d(\instruction_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_EX[17]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_EX[17] .is_wysiwyg = "true";
defparam \instruction_EX[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N9
dffeas \wsel_M[1] (
	.clk(CLK),
	.d(\wsel_M~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(wsel_M[1]),
	.prn(vcc));
// synopsys translate_off
defparam \wsel_M[1] .is_wysiwyg = "true";
defparam \wsel_M[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N3
dffeas \wsel_M[0] (
	.clk(CLK),
	.d(\wsel_M~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(wsel_M[0]),
	.prn(vcc));
// synopsys translate_off
defparam \wsel_M[0] .is_wysiwyg = "true";
defparam \wsel_M[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N15
dffeas \instruction_EX[18] (
	.clk(CLK),
	.d(\instruction_EX~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_EX[18]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_EX[18] .is_wysiwyg = "true";
defparam \instruction_EX[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N25
dffeas \instruction_EX[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instruction_EX~3_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_EX[19]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_EX[19] .is_wysiwyg = "true";
defparam \instruction_EX[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N27
dffeas \wsel_M[3] (
	.clk(CLK),
	.d(\wsel_M~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(wsel_M[3]),
	.prn(vcc));
// synopsys translate_off
defparam \wsel_M[3] .is_wysiwyg = "true";
defparam \wsel_M[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N5
dffeas \wsel_M[2] (
	.clk(CLK),
	.d(\wsel_M~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(wsel_M[2]),
	.prn(vcc));
// synopsys translate_off
defparam \wsel_M[2] .is_wysiwyg = "true";
defparam \wsel_M[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N25
dffeas \instruction_EX[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instruction_EX~4_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_EX[20]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_EX[20] .is_wysiwyg = "true";
defparam \instruction_EX[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y35_N21
dffeas \wsel_M[4] (
	.clk(CLK),
	.d(\wsel_M~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(wsel_M[4]),
	.prn(vcc));
// synopsys translate_off
defparam \wsel_M[4] .is_wysiwyg = "true";
defparam \wsel_M[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N7
dffeas \instruction_EX[22] (
	.clk(CLK),
	.d(\instruction_EX~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_EX[22]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_EX[22] .is_wysiwyg = "true";
defparam \instruction_EX[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N1
dffeas \instruction_EX[24] (
	.clk(CLK),
	.d(\instruction_EX~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_EX[24]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_EX[24] .is_wysiwyg = "true";
defparam \instruction_EX[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N19
dffeas \instruction_EX[23] (
	.clk(CLK),
	.d(\instruction_EX~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_EX[23]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_EX[23] .is_wysiwyg = "true";
defparam \instruction_EX[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N25
dffeas \instruction_EX[25] (
	.clk(CLK),
	.d(\instruction_EX~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_EX[25]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_EX[25] .is_wysiwyg = "true";
defparam \instruction_EX[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N1
dffeas \wsel_WB[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(wsel_M[1]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(wsel_WB[1]),
	.prn(vcc));
// synopsys translate_off
defparam \wsel_WB[1] .is_wysiwyg = "true";
defparam \wsel_WB[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N23
dffeas \wsel_WB[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(wsel_M[0]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(wsel_WB[0]),
	.prn(vcc));
// synopsys translate_off
defparam \wsel_WB[0] .is_wysiwyg = "true";
defparam \wsel_WB[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N13
dffeas \wsel_WB[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(wsel_M[3]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(wsel_WB[3]),
	.prn(vcc));
// synopsys translate_off
defparam \wsel_WB[3] .is_wysiwyg = "true";
defparam \wsel_WB[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N15
dffeas \wsel_WB[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(wsel_M[2]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(wsel_WB[2]),
	.prn(vcc));
// synopsys translate_off
defparam \wsel_WB[2] .is_wysiwyg = "true";
defparam \wsel_WB[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N3
dffeas \wsel_WB[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(wsel_M[4]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(wsel_WB[4]),
	.prn(vcc));
// synopsys translate_off
defparam \wsel_WB[4] .is_wysiwyg = "true";
defparam \wsel_WB[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N13
dffeas \ALUOp_EX[0] (
	.clk(CLK),
	.d(\ALUOp_EX~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUOp_EX[0]),
	.prn(vcc));
// synopsys translate_off
defparam \ALUOp_EX[0] .is_wysiwyg = "true";
defparam \ALUOp_EX[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N19
dffeas \ALUOp_EX[1] (
	.clk(CLK),
	.d(\ALUOp_EX~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUOp_EX[1]),
	.prn(vcc));
// synopsys translate_off
defparam \ALUOp_EX[1] .is_wysiwyg = "true";
defparam \ALUOp_EX[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N23
dffeas \ALUOp_EX[2] (
	.clk(CLK),
	.d(\ALUOp_EX~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUOp_EX[2]),
	.prn(vcc));
// synopsys translate_off
defparam \ALUOp_EX[2] .is_wysiwyg = "true";
defparam \ALUOp_EX[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N13
dffeas \ALUOp_EX[3] (
	.clk(CLK),
	.d(\ALUOp_EX~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ALUOp_EX[3]),
	.prn(vcc));
// synopsys translate_off
defparam \ALUOp_EX[3] .is_wysiwyg = "true";
defparam \ALUOp_EX[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N25
dffeas beq_EX(
	.clk(CLK),
	.d(\beq_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\beq_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam beq_EX.is_wysiwyg = "true";
defparam beq_EX.power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N31
dffeas bne_EX(
	.clk(CLK),
	.d(\bne_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bne_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam bne_EX.is_wysiwyg = "true";
defparam bne_EX.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N31
dffeas ALUSrc_EX(
	.clk(CLK),
	.d(\ALUSrc_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\ALUSrc_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam ALUSrc_EX.is_wysiwyg = "true";
defparam ALUSrc_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N20
cycloneive_lcell_comb \portB~15 (
// Equation(s):
// \portB~15_combout  = (\portB~14_combout  & (((\Equal3~2_combout )))) # (!\portB~14_combout  & ((\Equal3~2_combout  & (\wdat_WB[31]~3_combout )) # (!\Equal3~2_combout  & ((rdata2_EX[31])))))

	.dataa(\wdat_WB[31]~3_combout ),
	.datab(rdata2_EX[31]),
	.datac(\portB~14_combout ),
	.datad(\Equal3~2_combout ),
	.cin(gnd),
	.combout(\portB~15_combout ),
	.cout());
// synopsys translate_off
defparam \portB~15 .lut_mask = 16'hFA0C;
defparam \portB~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N22
cycloneive_lcell_comb \portB~16 (
// Equation(s):
// \portB~16_combout  = (\portB~14_combout  & ((\portB~15_combout  & ((\sw_forwarding_output~0_combout ))) # (!\portB~15_combout  & (\sign_ext[16]~0_combout )))) # (!\portB~14_combout  & (((\portB~15_combout ))))

	.dataa(\portB~14_combout ),
	.datab(\sign_ext[16]~0_combout ),
	.datac(\sw_forwarding_output~0_combout ),
	.datad(\portB~15_combout ),
	.cin(gnd),
	.combout(\portB~16_combout ),
	.cout());
// synopsys translate_off
defparam \portB~16 .lut_mask = 16'hF588;
defparam \portB~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N4
cycloneive_lcell_comb \portB~17 (
// Equation(s):
// \portB~17_combout  = (\portB~16_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(\ShiftOp_EX~q ),
	.datab(gnd),
	.datac(\portB~16_combout ),
	.datad(\Equal3~2_combout ),
	.cin(gnd),
	.combout(\portB~17_combout ),
	.cout());
// synopsys translate_off
defparam \portB~17 .lut_mask = 16'hF050;
defparam \portB~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N11
dffeas \dmemload_WB[30] (
	.clk(CLK),
	.d(\dpif.dmemload [30]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[30]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[30] .is_wysiwyg = "true";
defparam \dmemload_WB[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N23
dffeas \dmemload_WB[28] (
	.clk(CLK),
	.d(\dpif.dmemload [28]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[28]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[28] .is_wysiwyg = "true";
defparam \dmemload_WB[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N13
dffeas \pc_plus_4_WB[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[28]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[28]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[28] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N21
dffeas \dmemload_WB[27] (
	.clk(CLK),
	.d(\dpif.dmemload [27]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[27]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[27] .is_wysiwyg = "true";
defparam \dmemload_WB[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N31
dffeas \imm_WB[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[11]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[11]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[11] .is_wysiwyg = "true";
defparam \imm_WB[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N0
cycloneive_lcell_comb \portB~27 (
// Equation(s):
// \portB~27_combout  = (\portB~14_combout  & (((\Equal3~2_combout )))) # (!\portB~14_combout  & ((\Equal3~2_combout  & ((\wdat_WB[27]~11_combout ))) # (!\Equal3~2_combout  & (rdata2_EX[27]))))

	.dataa(rdata2_EX[27]),
	.datab(\wdat_WB[27]~11_combout ),
	.datac(\portB~14_combout ),
	.datad(\Equal3~2_combout ),
	.cin(gnd),
	.combout(\portB~27_combout ),
	.cout());
// synopsys translate_off
defparam \portB~27 .lut_mask = 16'hFC0A;
defparam \portB~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N24
cycloneive_lcell_comb \portB~28 (
// Equation(s):
// \portB~28_combout  = (\portB~14_combout  & ((\portB~27_combout  & (\sw_forwarding_output~4_combout )) # (!\portB~27_combout  & ((\sign_ext[16]~0_combout ))))) # (!\portB~14_combout  & (((\portB~27_combout ))))

	.dataa(\sw_forwarding_output~4_combout ),
	.datab(\sign_ext[16]~0_combout ),
	.datac(\portB~14_combout ),
	.datad(\portB~27_combout ),
	.cin(gnd),
	.combout(\portB~28_combout ),
	.cout());
// synopsys translate_off
defparam \portB~28 .lut_mask = 16'hAFC0;
defparam \portB~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N30
cycloneive_lcell_comb \portB~29 (
// Equation(s):
// \portB~29_combout  = (\portB~28_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(\Equal3~2_combout ),
	.datab(\ShiftOp_EX~q ),
	.datac(gnd),
	.datad(\portB~28_combout ),
	.cin(gnd),
	.combout(\portB~29_combout ),
	.cout());
// synopsys translate_off
defparam \portB~29 .lut_mask = 16'hBB00;
defparam \portB~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N8
cycloneive_lcell_comb \sw_forwarding_output~5 (
// Equation(s):
// \sw_forwarding_output~5_combout  = (\lui_M~q  & (imm_M[10])) # (!\lui_M~q  & ((porto_M_26)))

	.dataa(\lui_M~q ),
	.datab(imm_M[10]),
	.datac(porto_M_26),
	.datad(gnd),
	.cin(gnd),
	.combout(\sw_forwarding_output~5_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~5 .lut_mask = 16'hD8D8;
defparam \sw_forwarding_output~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N14
cycloneive_lcell_comb \portB~33 (
// Equation(s):
// \portB~33_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & (\sign_ext[16]~0_combout )) # (!\portB~14_combout  & ((rdata2_EX[25])))))

	.dataa(\portB~14_combout ),
	.datab(\ShiftOp_EX~q ),
	.datac(\sign_ext[16]~0_combout ),
	.datad(rdata2_EX[25]),
	.cin(gnd),
	.combout(\portB~33_combout ),
	.cout());
// synopsys translate_off
defparam \portB~33 .lut_mask = 16'h3120;
defparam \portB~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N20
cycloneive_lcell_comb \portB~34 (
// Equation(s):
// \portB~34_combout  = (\portB~14_combout  & ((\sw_forwarding_output~6_combout ))) # (!\portB~14_combout  & (\wdat_WB[25]~15_combout ))

	.dataa(\portB~14_combout ),
	.datab(\wdat_WB[25]~15_combout ),
	.datac(\sw_forwarding_output~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\portB~34_combout ),
	.cout());
// synopsys translate_off
defparam \portB~34 .lut_mask = 16'hE4E4;
defparam \portB~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N10
cycloneive_lcell_comb \portB~35 (
// Equation(s):
// \portB~35_combout  = (\Equal3~2_combout  & ((\portB~34_combout ))) # (!\Equal3~2_combout  & (\portB~33_combout ))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~33_combout ),
	.datad(\portB~34_combout ),
	.cin(gnd),
	.combout(\portB~35_combout ),
	.cout());
// synopsys translate_off
defparam \portB~35 .lut_mask = 16'hFA50;
defparam \portB~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N12
cycloneive_lcell_comb \portB~36 (
// Equation(s):
// \portB~36_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & ((\sign_ext[16]~0_combout ))) # (!\portB~14_combout  & (rdata2_EX[24]))))

	.dataa(\portB~14_combout ),
	.datab(rdata2_EX[24]),
	.datac(\sign_ext[16]~0_combout ),
	.datad(\ShiftOp_EX~q ),
	.cin(gnd),
	.combout(\portB~36_combout ),
	.cout());
// synopsys translate_off
defparam \portB~36 .lut_mask = 16'h00E4;
defparam \portB~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N8
cycloneive_lcell_comb \portB~37 (
// Equation(s):
// \portB~37_combout  = (\portB~14_combout  & (\sw_forwarding_output~7_combout )) # (!\portB~14_combout  & ((\wdat_WB[24]~17_combout )))

	.dataa(\portB~14_combout ),
	.datab(\sw_forwarding_output~7_combout ),
	.datac(\wdat_WB[24]~17_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\portB~37_combout ),
	.cout());
// synopsys translate_off
defparam \portB~37 .lut_mask = 16'hD8D8;
defparam \portB~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N6
cycloneive_lcell_comb \portB~38 (
// Equation(s):
// \portB~38_combout  = (\Equal3~2_combout  & (\portB~37_combout )) # (!\Equal3~2_combout  & ((\portB~36_combout )))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~37_combout ),
	.datad(\portB~36_combout ),
	.cin(gnd),
	.combout(\portB~38_combout ),
	.cout());
// synopsys translate_off
defparam \portB~38 .lut_mask = 16'hF5A0;
defparam \portB~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N30
cycloneive_lcell_comb \portB~39 (
// Equation(s):
// \portB~39_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & ((\sign_ext[16]~0_combout ))) # (!\portB~14_combout  & (rdata2_EX[23]))))

	.dataa(rdata2_EX[23]),
	.datab(\ShiftOp_EX~q ),
	.datac(\sign_ext[16]~0_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~39_combout ),
	.cout());
// synopsys translate_off
defparam \portB~39 .lut_mask = 16'h3022;
defparam \portB~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N0
cycloneive_lcell_comb \portB~40 (
// Equation(s):
// \portB~40_combout  = (\portB~14_combout  & (\sw_forwarding_output~8_combout )) # (!\portB~14_combout  & ((\wdat_WB[23]~19_combout )))

	.dataa(gnd),
	.datab(\sw_forwarding_output~8_combout ),
	.datac(\portB~14_combout ),
	.datad(\wdat_WB[23]~19_combout ),
	.cin(gnd),
	.combout(\portB~40_combout ),
	.cout());
// synopsys translate_off
defparam \portB~40 .lut_mask = 16'hCFC0;
defparam \portB~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N10
cycloneive_lcell_comb \portB~41 (
// Equation(s):
// \portB~41_combout  = (\Equal3~2_combout  & ((\portB~40_combout ))) # (!\Equal3~2_combout  & (\portB~39_combout ))

	.dataa(gnd),
	.datab(\Equal3~2_combout ),
	.datac(\portB~39_combout ),
	.datad(\portB~40_combout ),
	.cin(gnd),
	.combout(\portB~41_combout ),
	.cout());
// synopsys translate_off
defparam \portB~41 .lut_mask = 16'hFC30;
defparam \portB~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N16
cycloneive_lcell_comb \portB~42 (
// Equation(s):
// \portB~42_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & ((\sign_ext[16]~0_combout ))) # (!\portB~14_combout  & (rdata2_EX[22]))))

	.dataa(rdata2_EX[22]),
	.datab(\ShiftOp_EX~q ),
	.datac(\portB~14_combout ),
	.datad(\sign_ext[16]~0_combout ),
	.cin(gnd),
	.combout(\portB~42_combout ),
	.cout());
// synopsys translate_off
defparam \portB~42 .lut_mask = 16'h3202;
defparam \portB~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N30
cycloneive_lcell_comb \sw_forwarding_output~9 (
// Equation(s):
// \sw_forwarding_output~9_combout  = (\lui_M~q  & (imm_M[6])) # (!\lui_M~q  & ((porto_M_22)))

	.dataa(gnd),
	.datab(imm_M[6]),
	.datac(\lui_M~q ),
	.datad(porto_M_22),
	.cin(gnd),
	.combout(\sw_forwarding_output~9_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~9 .lut_mask = 16'hCFC0;
defparam \sw_forwarding_output~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N22
cycloneive_lcell_comb \portB~43 (
// Equation(s):
// \portB~43_combout  = (\portB~14_combout  & (\sw_forwarding_output~9_combout )) # (!\portB~14_combout  & ((\wdat_WB[22]~21_combout )))

	.dataa(\sw_forwarding_output~9_combout ),
	.datab(gnd),
	.datac(\portB~14_combout ),
	.datad(\wdat_WB[22]~21_combout ),
	.cin(gnd),
	.combout(\portB~43_combout ),
	.cout());
// synopsys translate_off
defparam \portB~43 .lut_mask = 16'hAFA0;
defparam \portB~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N12
cycloneive_lcell_comb \portB~44 (
// Equation(s):
// \portB~44_combout  = (\Equal3~2_combout  & (\portB~43_combout )) # (!\Equal3~2_combout  & ((\portB~42_combout )))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~43_combout ),
	.datad(\portB~42_combout ),
	.cin(gnd),
	.combout(\portB~44_combout ),
	.cout());
// synopsys translate_off
defparam \portB~44 .lut_mask = 16'hF5A0;
defparam \portB~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N15
dffeas \pc_plus_4_WB[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[21]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[21]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[21] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N11
dffeas \dmemload_WB[21] (
	.clk(CLK),
	.d(\dpif.dmemload [21]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[21]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[21] .is_wysiwyg = "true";
defparam \dmemload_WB[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N2
cycloneive_lcell_comb \portB~48 (
// Equation(s):
// \portB~48_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & (\sign_ext[16]~0_combout )) # (!\portB~14_combout  & ((rdata2_EX[20])))))

	.dataa(\portB~14_combout ),
	.datab(\ShiftOp_EX~q ),
	.datac(\sign_ext[16]~0_combout ),
	.datad(rdata2_EX[20]),
	.cin(gnd),
	.combout(\portB~48_combout ),
	.cout());
// synopsys translate_off
defparam \portB~48 .lut_mask = 16'h3120;
defparam \portB~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N8
cycloneive_lcell_comb \portB~49 (
// Equation(s):
// \portB~49_combout  = (\portB~14_combout  & ((\sw_forwarding_output~11_combout ))) # (!\portB~14_combout  & (\wdat_WB[20]~25_combout ))

	.dataa(\wdat_WB[20]~25_combout ),
	.datab(\sw_forwarding_output~11_combout ),
	.datac(\portB~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\portB~49_combout ),
	.cout());
// synopsys translate_off
defparam \portB~49 .lut_mask = 16'hCACA;
defparam \portB~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N6
cycloneive_lcell_comb \portB~50 (
// Equation(s):
// \portB~50_combout  = (\Equal3~2_combout  & (\portB~49_combout )) # (!\Equal3~2_combout  & ((\portB~48_combout )))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~49_combout ),
	.datad(\portB~48_combout ),
	.cin(gnd),
	.combout(\portB~50_combout ),
	.cout());
// synopsys translate_off
defparam \portB~50 .lut_mask = 16'hF5A0;
defparam \portB~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N23
dffeas \dmemload_WB[19] (
	.clk(CLK),
	.d(\dmemload_WB[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[19]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[19] .is_wysiwyg = "true";
defparam \dmemload_WB[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N31
dffeas \dmemload_WB[18] (
	.clk(CLK),
	.d(\dmemload_WB[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[18]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[18] .is_wysiwyg = "true";
defparam \dmemload_WB[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N13
dffeas \pc_plus_4_WB[18] (
	.clk(CLK),
	.d(\pc_plus_4_WB[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[18]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[18] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N28
cycloneive_lcell_comb \portB~57 (
// Equation(s):
// \portB~57_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & ((\sign_ext[16]~0_combout ))) # (!\portB~14_combout  & (rdata2_EX[17]))))

	.dataa(\ShiftOp_EX~q ),
	.datab(rdata2_EX[17]),
	.datac(\sign_ext[16]~0_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~57_combout ),
	.cout());
// synopsys translate_off
defparam \portB~57 .lut_mask = 16'h5044;
defparam \portB~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y28_N9
dffeas \dmemload_WB[17] (
	.clk(CLK),
	.d(\dpif.dmemload [17]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[17]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[17] .is_wysiwyg = "true";
defparam \dmemload_WB[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N27
dffeas \imm_WB[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[1]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[1]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[1] .is_wysiwyg = "true";
defparam \imm_WB[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N4
cycloneive_lcell_comb \portB~58 (
// Equation(s):
// \portB~58_combout  = (\portB~14_combout  & ((\sw_forwarding_output~14_combout ))) # (!\portB~14_combout  & (\wdat_WB[17]~31_combout ))

	.dataa(\wdat_WB[17]~31_combout ),
	.datab(\sw_forwarding_output~14_combout ),
	.datac(gnd),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~58_combout ),
	.cout());
// synopsys translate_off
defparam \portB~58 .lut_mask = 16'hCCAA;
defparam \portB~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N22
cycloneive_lcell_comb \portB~59 (
// Equation(s):
// \portB~59_combout  = (\Equal3~2_combout  & (\portB~58_combout )) # (!\Equal3~2_combout  & ((\portB~57_combout )))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~58_combout ),
	.datad(\portB~57_combout ),
	.cin(gnd),
	.combout(\portB~59_combout ),
	.cout());
// synopsys translate_off
defparam \portB~59 .lut_mask = 16'hF5A0;
defparam \portB~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N12
cycloneive_lcell_comb \portB~60 (
// Equation(s):
// \portB~60_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & ((\sign_ext[16]~0_combout ))) # (!\portB~14_combout  & (rdata2_EX[16]))))

	.dataa(\ShiftOp_EX~q ),
	.datab(rdata2_EX[16]),
	.datac(\sign_ext[16]~0_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~60_combout ),
	.cout());
// synopsys translate_off
defparam \portB~60 .lut_mask = 16'h5044;
defparam \portB~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N23
dffeas \pc_plus_4_WB[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[16]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[16]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[16] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N1
dffeas \dmemload_WB[15] (
	.clk(CLK),
	.d(\dmemload_WB[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[15]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[15] .is_wysiwyg = "true";
defparam \dmemload_WB[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N23
dffeas \dmemload_WB[14] (
	.clk(CLK),
	.d(\dpif.dmemload [14]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[14]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[14] .is_wysiwyg = "true";
defparam \dmemload_WB[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N16
cycloneive_lcell_comb \sw_forwarding_output~17 (
// Equation(s):
// \sw_forwarding_output~17_combout  = (!\lui_M~q  & porto_M_14)

	.dataa(\lui_M~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(porto_M_14),
	.cin(gnd),
	.combout(\sw_forwarding_output~17_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~17 .lut_mask = 16'h5500;
defparam \sw_forwarding_output~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N4
cycloneive_lcell_comb \portB~67 (
// Equation(s):
// \portB~67_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & ((imm_EX[13]))) # (!\portB~14_combout  & (rdata2_EX[13]))))

	.dataa(rdata2_EX[13]),
	.datab(imm_EX[13]),
	.datac(\ShiftOp_EX~q ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~67_combout ),
	.cout());
// synopsys translate_off
defparam \portB~67 .lut_mask = 16'h0C0A;
defparam \portB~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N30
cycloneive_lcell_comb \portB~68 (
// Equation(s):
// \portB~68_combout  = (\Equal3~2_combout  & ((\portB~112_combout ))) # (!\Equal3~2_combout  & (\portB~67_combout ))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~67_combout ),
	.datad(\portB~112_combout ),
	.cin(gnd),
	.combout(\portB~68_combout ),
	.cout());
// synopsys translate_off
defparam \portB~68 .lut_mask = 16'hFA50;
defparam \portB~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N8
cycloneive_lcell_comb \portB~69 (
// Equation(s):
// \portB~69_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & ((imm_EX[12]))) # (!\portB~14_combout  & (rdata2_EX[12]))))

	.dataa(rdata2_EX[12]),
	.datab(imm_EX[12]),
	.datac(\ShiftOp_EX~q ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~69_combout ),
	.cout());
// synopsys translate_off
defparam \portB~69 .lut_mask = 16'h0C0A;
defparam \portB~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N26
cycloneive_lcell_comb \portB~70 (
// Equation(s):
// \portB~70_combout  = (\Equal3~2_combout  & ((\portB~113_combout ))) # (!\Equal3~2_combout  & (\portB~69_combout ))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~69_combout ),
	.datad(\portB~113_combout ),
	.cin(gnd),
	.combout(\portB~70_combout ),
	.cout());
// synopsys translate_off
defparam \portB~70 .lut_mask = 16'hFA50;
defparam \portB~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N13
dffeas \dmemload_WB[8] (
	.clk(CLK),
	.d(\dpif.dmemload [8]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[8]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[8] .is_wysiwyg = "true";
defparam \dmemload_WB[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N16
cycloneive_lcell_comb \portB~74 (
// Equation(s):
// \portB~74_combout  = (\Equal3~2_combout  & ((\sw_forwarding_output~21_combout ) # ((!\portB~14_combout )))) # (!\Equal3~2_combout  & (((imm_EX[8] & \portB~14_combout ))))

	.dataa(\sw_forwarding_output~21_combout ),
	.datab(imm_EX[8]),
	.datac(\Equal3~2_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~74_combout ),
	.cout());
// synopsys translate_off
defparam \portB~74 .lut_mask = 16'hACF0;
defparam \portB~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N26
cycloneive_lcell_comb \portB~75 (
// Equation(s):
// \portB~75_combout  = (\portB~14_combout  & (((\portB~74_combout )))) # (!\portB~14_combout  & ((\portB~74_combout  & (\wdat_WB[8]~45_combout )) # (!\portB~74_combout  & ((rdata2_EX[8])))))

	.dataa(\wdat_WB[8]~45_combout ),
	.datab(rdata2_EX[8]),
	.datac(\portB~14_combout ),
	.datad(\portB~74_combout ),
	.cin(gnd),
	.combout(\portB~75_combout ),
	.cout());
// synopsys translate_off
defparam \portB~75 .lut_mask = 16'hFA0C;
defparam \portB~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N28
cycloneive_lcell_comb \portB~76 (
// Equation(s):
// \portB~76_combout  = (\portB~75_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~75_combout ),
	.datad(\ShiftOp_EX~q ),
	.cin(gnd),
	.combout(\portB~76_combout ),
	.cout());
// synopsys translate_off
defparam \portB~76 .lut_mask = 16'hA0F0;
defparam \portB~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N29
dffeas \imm_EX[11] (
	.clk(CLK),
	.d(\imm_EX~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[11]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[11] .is_wysiwyg = "true";
defparam \imm_EX[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N25
dffeas \dmemload_WB[11] (
	.clk(CLK),
	.d(\dpif.dmemload [11]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[11]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[11] .is_wysiwyg = "true";
defparam \dmemload_WB[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N6
cycloneive_lcell_comb \portB~77 (
// Equation(s):
// \portB~77_combout  = (\Equal3~2_combout  & ((\wdat_WB[11]~47_combout ) # ((\portB~14_combout )))) # (!\Equal3~2_combout  & (((rdata2_EX[11] & !\portB~14_combout ))))

	.dataa(\wdat_WB[11]~47_combout ),
	.datab(rdata2_EX[11]),
	.datac(\Equal3~2_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~77_combout ),
	.cout());
// synopsys translate_off
defparam \portB~77 .lut_mask = 16'hF0AC;
defparam \portB~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N0
cycloneive_lcell_comb \portB~78 (
// Equation(s):
// \portB~78_combout  = (\portB~14_combout  & ((\portB~77_combout  & (\sw_forwarding_output~22_combout )) # (!\portB~77_combout  & ((imm_EX[11]))))) # (!\portB~14_combout  & (((\portB~77_combout ))))

	.dataa(\sw_forwarding_output~22_combout ),
	.datab(imm_EX[11]),
	.datac(\portB~14_combout ),
	.datad(\portB~77_combout ),
	.cin(gnd),
	.combout(\portB~78_combout ),
	.cout());
// synopsys translate_off
defparam \portB~78 .lut_mask = 16'hAFC0;
defparam \portB~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N11
dffeas \dmemload_WB[10] (
	.clk(CLK),
	.d(\dpif.dmemload [10]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[10]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[10] .is_wysiwyg = "true";
defparam \dmemload_WB[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N18
cycloneive_lcell_comb \portB~79 (
// Equation(s):
// \portB~79_combout  = (\Equal3~2_combout  & (((\portB~14_combout )))) # (!\Equal3~2_combout  & ((\portB~14_combout  & (imm_EX[10])) # (!\portB~14_combout  & ((rdata2_EX[10])))))

	.dataa(imm_EX[10]),
	.datab(rdata2_EX[10]),
	.datac(\Equal3~2_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~79_combout ),
	.cout());
// synopsys translate_off
defparam \portB~79 .lut_mask = 16'hFA0C;
defparam \portB~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N12
cycloneive_lcell_comb \portB~80 (
// Equation(s):
// \portB~80_combout  = (\Equal3~2_combout  & ((\portB~79_combout  & (\sw_forwarding_output~23_combout )) # (!\portB~79_combout  & ((\wdat_WB[10]~49_combout ))))) # (!\Equal3~2_combout  & (((\portB~79_combout ))))

	.dataa(\sw_forwarding_output~23_combout ),
	.datab(\wdat_WB[10]~49_combout ),
	.datac(\Equal3~2_combout ),
	.datad(\portB~79_combout ),
	.cin(gnd),
	.combout(\portB~80_combout ),
	.cout());
// synopsys translate_off
defparam \portB~80 .lut_mask = 16'hAFC0;
defparam \portB~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N4
cycloneive_lcell_comb \portB~81 (
// Equation(s):
// \portB~81_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & ((imm_EX[7]))) # (!\portB~14_combout  & (rdata2_EX[7]))))

	.dataa(rdata2_EX[7]),
	.datab(\ShiftOp_EX~q ),
	.datac(imm_EX[7]),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~81_combout ),
	.cout());
// synopsys translate_off
defparam \portB~81 .lut_mask = 16'h3022;
defparam \portB~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N30
cycloneive_lcell_comb \portB~82 (
// Equation(s):
// \portB~82_combout  = (\Equal3~2_combout  & ((\portB~114_combout ))) # (!\Equal3~2_combout  & (\portB~81_combout ))

	.dataa(gnd),
	.datab(\portB~81_combout ),
	.datac(\portB~114_combout ),
	.datad(\Equal3~2_combout ),
	.cin(gnd),
	.combout(\portB~82_combout ),
	.cout());
// synopsys translate_off
defparam \portB~82 .lut_mask = 16'hF0CC;
defparam \portB~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N27
dffeas \dmemload_WB[6] (
	.clk(CLK),
	.d(\dpif.dmemload [6]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[6]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[6] .is_wysiwyg = "true";
defparam \dmemload_WB[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N0
cycloneive_lcell_comb \sw_forwarding_output~25 (
// Equation(s):
// \sw_forwarding_output~25_combout  = (!\lui_M~q  & porto_M_6)

	.dataa(\lui_M~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(porto_M_6),
	.cin(gnd),
	.combout(\sw_forwarding_output~25_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~25 .lut_mask = 16'h5500;
defparam \sw_forwarding_output~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N4
cycloneive_lcell_comb \portB~85 (
// Equation(s):
// \portB~85_combout  = (\ALUSrc_EX~q  & ((imm_EX[5]))) # (!\ALUSrc_EX~q  & (rdata2_EX[5]))

	.dataa(\ALUSrc_EX~q ),
	.datab(rdata2_EX[5]),
	.datac(imm_EX[5]),
	.datad(gnd),
	.cin(gnd),
	.combout(\portB~85_combout ),
	.cout());
// synopsys translate_off
defparam \portB~85 .lut_mask = 16'hE4E4;
defparam \portB~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N2
cycloneive_lcell_comb \portB~86 (
// Equation(s):
// \portB~86_combout  = (fuifforward_B_11 & ((\wdat_WB[5]~55_combout ))) # (!fuifforward_B_11 & (\portB~85_combout ))

	.dataa(gnd),
	.datab(\portB~85_combout ),
	.datac(\wdat_WB[5]~55_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_B[1]~4_combout ),
	.cin(gnd),
	.combout(\portB~86_combout ),
	.cout());
// synopsys translate_off
defparam \portB~86 .lut_mask = 16'hF0CC;
defparam \portB~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N24
cycloneive_lcell_comb \portB~87 (
// Equation(s):
// \portB~87_combout  = (\portB~116_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(gnd),
	.datab(\ShiftOp_EX~q ),
	.datac(\Equal3~2_combout ),
	.datad(\portB~116_combout ),
	.cin(gnd),
	.combout(\portB~87_combout ),
	.cout());
// synopsys translate_off
defparam \portB~87 .lut_mask = 16'hF300;
defparam \portB~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N26
cycloneive_lcell_comb \portA~8 (
// Equation(s):
// \portA~8_combout  = (fuifforward_A_01 & (porto_M_2 & ((!\lui_M~q )))) # (!fuifforward_A_01 & (((rdata1_EX[2]))))

	.dataa(porto_M_2),
	.datab(rdata1_EX[2]),
	.datac(\lui_M~q ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~8_combout ),
	.cout());
// synopsys translate_off
defparam \portA~8 .lut_mask = 16'h0ACC;
defparam \portA~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N28
cycloneive_lcell_comb \portA~9 (
// Equation(s):
// \portA~9_combout  = (fuifforward_A_11 & (\wdat_WB[2]~57_combout )) # (!fuifforward_A_11 & ((\portA~8_combout )))

	.dataa(\wdat_WB[2]~57_combout ),
	.datab(gnd),
	.datac(\portA~8_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.cin(gnd),
	.combout(\portA~9_combout ),
	.cout());
// synopsys translate_off
defparam \portA~9 .lut_mask = 16'hAAF0;
defparam \portA~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N16
cycloneive_lcell_comb \portA~10 (
// Equation(s):
// \portA~10_combout  = (\regWrite_M~q  & (fuifforward_A_0 & ((instruction_EX[21]) # (!Equal3))))

	.dataa(\regWrite_M~q ),
	.datab(instruction_EX[21]),
	.datac(\FORWARDING_UNIT|Equal3~0_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~2_combout ),
	.cin(gnd),
	.combout(\portA~10_combout ),
	.cout());
// synopsys translate_off
defparam \portA~10 .lut_mask = 16'h8A00;
defparam \portA~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N10
cycloneive_lcell_comb \portA~11 (
// Equation(s):
// \portA~11_combout  = (\portA~10_combout  & (((porto_M_1 & !\lui_M~q )))) # (!\portA~10_combout  & (rdata1_EX[1]))

	.dataa(rdata1_EX[1]),
	.datab(porto_M_1),
	.datac(\lui_M~q ),
	.datad(\portA~10_combout ),
	.cin(gnd),
	.combout(\portA~11_combout ),
	.cout());
// synopsys translate_off
defparam \portA~11 .lut_mask = 16'h0CAA;
defparam \portA~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N20
cycloneive_lcell_comb \portA~12 (
// Equation(s):
// \portA~12_combout  = (fuifforward_A_11 & (\wdat_WB[1]~59_combout )) # (!fuifforward_A_11 & ((\portA~11_combout )))

	.dataa(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datab(gnd),
	.datac(\wdat_WB[1]~59_combout ),
	.datad(\portA~11_combout ),
	.cin(gnd),
	.combout(\portA~12_combout ),
	.cout());
// synopsys translate_off
defparam \portA~12 .lut_mask = 16'hF5A0;
defparam \portA~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N20
cycloneive_lcell_comb \portB~89 (
// Equation(s):
// \portB~89_combout  = (\ShiftOp_EX~q ) # ((!\ALUSrc_EX~q  & rdata2_EX[0]))

	.dataa(\ShiftOp_EX~q ),
	.datab(gnd),
	.datac(\ALUSrc_EX~q ),
	.datad(rdata2_EX[0]),
	.cin(gnd),
	.combout(\portB~89_combout ),
	.cout());
// synopsys translate_off
defparam \portB~89 .lut_mask = 16'hAFAA;
defparam \portB~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N22
cycloneive_lcell_comb \portB~90 (
// Equation(s):
// \portB~90_combout  = (\Equal2~0_combout  & (((\wdat_WB[0]~61_combout )))) # (!\Equal2~0_combout  & ((fuifforward_B_11 & ((\wdat_WB[0]~61_combout ))) # (!fuifforward_B_11 & (\portB~89_combout ))))

	.dataa(\Equal2~0_combout ),
	.datab(\portB~89_combout ),
	.datac(\wdat_WB[0]~61_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_B[1]~4_combout ),
	.cin(gnd),
	.combout(\portB~90_combout ),
	.cout());
// synopsys translate_off
defparam \portB~90 .lut_mask = 16'hF0E4;
defparam \portB~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N28
cycloneive_lcell_comb \portB~91 (
// Equation(s):
// \portB~91_combout  = (\portB~90_combout  & (((imm_EX[6]) # (!\portB~88_combout )))) # (!\portB~90_combout  & (imm_EX[0] & ((\portB~88_combout ))))

	.dataa(imm_EX[0]),
	.datab(imm_EX[6]),
	.datac(\portB~90_combout ),
	.datad(\portB~88_combout ),
	.cin(gnd),
	.combout(\portB~91_combout ),
	.cout());
// synopsys translate_off
defparam \portB~91 .lut_mask = 16'hCAF0;
defparam \portB~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N18
cycloneive_lcell_comb \portB~92 (
// Equation(s):
// \portB~92_combout  = (\Equal2~0_combout  & (porto_M_0 & (!\lui_M~q ))) # (!\Equal2~0_combout  & (((\portB~91_combout ))))

	.dataa(\Equal2~0_combout ),
	.datab(porto_M_0),
	.datac(\lui_M~q ),
	.datad(\portB~91_combout ),
	.cin(gnd),
	.combout(\portB~92_combout ),
	.cout());
// synopsys translate_off
defparam \portB~92 .lut_mask = 16'h5D08;
defparam \portB~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N22
cycloneive_lcell_comb \portB~94 (
// Equation(s):
// \portB~94_combout  = (\ALUSrc_EX~q  & ((imm_EX[1]))) # (!\ALUSrc_EX~q  & (rdata2_EX[1]))

	.dataa(gnd),
	.datab(rdata2_EX[1]),
	.datac(imm_EX[1]),
	.datad(\ALUSrc_EX~q ),
	.cin(gnd),
	.combout(\portB~94_combout ),
	.cout());
// synopsys translate_off
defparam \portB~94 .lut_mask = 16'hF0CC;
defparam \portB~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N0
cycloneive_lcell_comb \portB~95 (
// Equation(s):
// \portB~95_combout  = (!\Equal2~0_combout  & (!fuifforward_B_11 & ((\ShiftOp_EX~q ) # (\portB~94_combout ))))

	.dataa(\Equal2~0_combout ),
	.datab(\ShiftOp_EX~q ),
	.datac(\portB~94_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_B[1]~4_combout ),
	.cin(gnd),
	.combout(\portB~95_combout ),
	.cout());
// synopsys translate_off
defparam \portB~95 .lut_mask = 16'h0054;
defparam \portB~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N6
cycloneive_lcell_comb \portB~96 (
// Equation(s):
// \portB~96_combout  = (\portB~93_combout  & ((\portB~95_combout  & (imm_EX[7])) # (!\portB~95_combout  & ((\wdat_WB[1]~59_combout ))))) # (!\portB~93_combout  & (((\portB~95_combout ))))

	.dataa(imm_EX[7]),
	.datab(\wdat_WB[1]~59_combout ),
	.datac(\portB~93_combout ),
	.datad(\portB~95_combout ),
	.cin(gnd),
	.combout(\portB~96_combout ),
	.cout());
// synopsys translate_off
defparam \portB~96 .lut_mask = 16'hAFC0;
defparam \portB~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N12
cycloneive_lcell_comb \portB~97 (
// Equation(s):
// \portB~97_combout  = (\Equal2~0_combout  & (!\lui_M~q  & (porto_M_1))) # (!\Equal2~0_combout  & (((\portB~96_combout ))))

	.dataa(\Equal2~0_combout ),
	.datab(\lui_M~q ),
	.datac(porto_M_1),
	.datad(\portB~96_combout ),
	.cin(gnd),
	.combout(\portB~97_combout ),
	.cout());
// synopsys translate_off
defparam \portB~97 .lut_mask = 16'h7520;
defparam \portB~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N5
dffeas \dmemload_WB[4] (
	.clk(CLK),
	.d(\dmemload_WB[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[4]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[4] .is_wysiwyg = "true";
defparam \dmemload_WB[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N23
dffeas \porto_WB[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_4),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[4]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[4] .is_wysiwyg = "true";
defparam \porto_WB[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N22
cycloneive_lcell_comb \wdat_WB[4]~62 (
// Equation(s):
// \wdat_WB[4]~62_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[4])) # (!\memToReg_WB~q  & ((porto_WB[4])))))

	.dataa(dmemload_WB[4]),
	.datab(\jal_WB~q ),
	.datac(porto_WB[4]),
	.datad(\memToReg_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[4]~62_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[4]~62 .lut_mask = 16'h2230;
defparam \wdat_WB[4]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N2
cycloneive_lcell_comb \portA~13 (
// Equation(s):
// \portA~13_combout  = (fuifforward_A_01 & (porto_M_4 & (!\lui_M~q ))) # (!fuifforward_A_01 & (((rdata1_EX[4]))))

	.dataa(porto_M_4),
	.datab(\lui_M~q ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(rdata1_EX[4]),
	.cin(gnd),
	.combout(\portA~13_combout ),
	.cout());
// synopsys translate_off
defparam \portA~13 .lut_mask = 16'h2F20;
defparam \portA~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N20
cycloneive_lcell_comb \portA~14 (
// Equation(s):
// \portA~14_combout  = (fuifforward_A_11 & (\wdat_WB[4]~63_combout )) # (!fuifforward_A_11 & ((\portA~13_combout )))

	.dataa(\wdat_WB[4]~63_combout ),
	.datab(gnd),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~13_combout ),
	.cin(gnd),
	.combout(\portA~14_combout ),
	.cout());
// synopsys translate_off
defparam \portA~14 .lut_mask = 16'hAFA0;
defparam \portA~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N23
dffeas \dmemload_WB[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_3),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[3]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[3] .is_wysiwyg = "true";
defparam \dmemload_WB[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N14
cycloneive_lcell_comb \portA~15 (
// Equation(s):
// \portA~15_combout  = (fuifforward_A_01 & (porto_M_3 & (!\lui_M~q ))) # (!fuifforward_A_01 & (((rdata1_EX[3]))))

	.dataa(porto_M_3),
	.datab(\lui_M~q ),
	.datac(rdata1_EX[3]),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~15_combout ),
	.cout());
// synopsys translate_off
defparam \portA~15 .lut_mask = 16'h22F0;
defparam \portA~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N24
cycloneive_lcell_comb \portA~16 (
// Equation(s):
// \portA~16_combout  = (fuifforward_A_11 & (\wdat_WB[3]~65_combout )) # (!fuifforward_A_11 & ((\portA~15_combout )))

	.dataa(\wdat_WB[3]~65_combout ),
	.datab(gnd),
	.datac(\portA~15_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.cin(gnd),
	.combout(\portA~16_combout ),
	.cout());
// synopsys translate_off
defparam \portA~16 .lut_mask = 16'hAAF0;
defparam \portA~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N22
cycloneive_lcell_comb \portA~17 (
// Equation(s):
// \portA~17_combout  = (fuifforward_A_11 & (\wdat_WB[8]~45_combout )) # (!fuifforward_A_11 & ((\portA~70_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[8]~45_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~70_combout ),
	.cin(gnd),
	.combout(\portA~17_combout ),
	.cout());
// synopsys translate_off
defparam \portA~17 .lut_mask = 16'hCFC0;
defparam \portA~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N20
cycloneive_lcell_comb \portA~18 (
// Equation(s):
// \portA~18_combout  = (fuifforward_A_01 & (((porto_M_7 & !\lui_M~q )))) # (!fuifforward_A_01 & (rdata1_EX[7]))

	.dataa(rdata1_EX[7]),
	.datab(porto_M_7),
	.datac(\lui_M~q ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~18_combout ),
	.cout());
// synopsys translate_off
defparam \portA~18 .lut_mask = 16'h0CAA;
defparam \portA~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N6
cycloneive_lcell_comb \portA~19 (
// Equation(s):
// \portA~19_combout  = (fuifforward_A_11 & (\wdat_WB[7]~51_combout )) # (!fuifforward_A_11 & ((\portA~18_combout )))

	.dataa(\wdat_WB[7]~51_combout ),
	.datab(gnd),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~18_combout ),
	.cin(gnd),
	.combout(\portA~19_combout ),
	.cout());
// synopsys translate_off
defparam \portA~19 .lut_mask = 16'hAFA0;
defparam \portA~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N2
cycloneive_lcell_comb \portA~20 (
// Equation(s):
// \portA~20_combout  = (fuifforward_A_01 & (((!\lui_M~q  & porto_M_6)))) # (!fuifforward_A_01 & (rdata1_EX[6]))

	.dataa(rdata1_EX[6]),
	.datab(\lui_M~q ),
	.datac(porto_M_6),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~20_combout ),
	.cout());
// synopsys translate_off
defparam \portA~20 .lut_mask = 16'h30AA;
defparam \portA~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N24
cycloneive_lcell_comb \portA~21 (
// Equation(s):
// \portA~21_combout  = (fuifforward_A_11 & (\wdat_WB[6]~53_combout )) # (!fuifforward_A_11 & ((\portA~20_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[6]~53_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~20_combout ),
	.cin(gnd),
	.combout(\portA~21_combout ),
	.cout());
// synopsys translate_off
defparam \portA~21 .lut_mask = 16'hCFC0;
defparam \portA~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N12
cycloneive_lcell_comb \portA~22 (
// Equation(s):
// \portA~22_combout  = (fuifforward_A_01 & (porto_M_5 & ((!\lui_M~q )))) # (!fuifforward_A_01 & (((rdata1_EX[5]))))

	.dataa(porto_M_5),
	.datab(rdata1_EX[5]),
	.datac(\lui_M~q ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~22_combout ),
	.cout());
// synopsys translate_off
defparam \portA~22 .lut_mask = 16'h0ACC;
defparam \portA~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N30
cycloneive_lcell_comb \portA~23 (
// Equation(s):
// \portA~23_combout  = (fuifforward_A_11 & (\wdat_WB[5]~55_combout )) # (!fuifforward_A_11 & ((\portA~22_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[5]~55_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~22_combout ),
	.cin(gnd),
	.combout(\portA~23_combout ),
	.cout());
// synopsys translate_off
defparam \portA~23 .lut_mask = 16'hCFC0;
defparam \portA~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N10
cycloneive_lcell_comb \portB~101 (
// Equation(s):
// \portB~101_combout  = (\portB~88_combout  & (((imm_EX[3]) # (\portB~93_combout )))) # (!\portB~88_combout  & (rdata2_EX[3] & ((!\portB~93_combout ))))

	.dataa(rdata2_EX[3]),
	.datab(imm_EX[3]),
	.datac(\portB~88_combout ),
	.datad(\portB~93_combout ),
	.cin(gnd),
	.combout(\portB~101_combout ),
	.cout());
// synopsys translate_off
defparam \portB~101 .lut_mask = 16'hF0CA;
defparam \portB~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N16
cycloneive_lcell_comb \portB~102 (
// Equation(s):
// \portB~102_combout  = (\portB~93_combout  & ((\portB~101_combout  & (imm_EX[9])) # (!\portB~101_combout  & ((\wdat_WB[3]~65_combout ))))) # (!\portB~93_combout  & (((\portB~101_combout ))))

	.dataa(imm_EX[9]),
	.datab(\portB~93_combout ),
	.datac(\wdat_WB[3]~65_combout ),
	.datad(\portB~101_combout ),
	.cin(gnd),
	.combout(\portB~102_combout ),
	.cout());
// synopsys translate_off
defparam \portB~102 .lut_mask = 16'hBBC0;
defparam \portB~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N2
cycloneive_lcell_comb \portB~103 (
// Equation(s):
// \portB~103_combout  = (\Equal2~0_combout  & (porto_M_3 & (!\lui_M~q ))) # (!\Equal2~0_combout  & (((\portB~102_combout ))))

	.dataa(porto_M_3),
	.datab(\lui_M~q ),
	.datac(\Equal2~0_combout ),
	.datad(\portB~102_combout ),
	.cin(gnd),
	.combout(\portB~103_combout ),
	.cout());
// synopsys translate_off
defparam \portB~103 .lut_mask = 16'h2F20;
defparam \portB~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N4
cycloneive_lcell_comb \portA~24 (
// Equation(s):
// \portA~24_combout  = (fuifforward_A_01 & ((\sw_forwarding_output~15_combout ))) # (!fuifforward_A_01 & (rdata1_EX[16]))

	.dataa(rdata1_EX[16]),
	.datab(gnd),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(\sw_forwarding_output~15_combout ),
	.cin(gnd),
	.combout(\portA~24_combout ),
	.cout());
// synopsys translate_off
defparam \portA~24 .lut_mask = 16'hFA0A;
defparam \portA~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N6
cycloneive_lcell_comb \portA~25 (
// Equation(s):
// \portA~25_combout  = (fuifforward_A_11 & (\wdat_WB[16]~33_combout )) # (!fuifforward_A_11 & ((\portA~24_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[16]~33_combout ),
	.datac(\portA~24_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.cin(gnd),
	.combout(\portA~25_combout ),
	.cout());
// synopsys translate_off
defparam \portA~25 .lut_mask = 16'hCCF0;
defparam \portA~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N8
cycloneive_lcell_comb \portA~26 (
// Equation(s):
// \portA~26_combout  = (fuifforward_A_01 & (porto_M_15 & (!\lui_M~q ))) # (!fuifforward_A_01 & (((rdata1_EX[15]))))

	.dataa(porto_M_15),
	.datab(\lui_M~q ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(rdata1_EX[15]),
	.cin(gnd),
	.combout(\portA~26_combout ),
	.cout());
// synopsys translate_off
defparam \portA~26 .lut_mask = 16'h2F20;
defparam \portA~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N30
cycloneive_lcell_comb \portA~27 (
// Equation(s):
// \portA~27_combout  = (fuifforward_A_11 & (\wdat_WB[15]~35_combout )) # (!fuifforward_A_11 & ((\portA~26_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[15]~35_combout ),
	.datac(\portA~26_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.cin(gnd),
	.combout(\portA~27_combout ),
	.cout());
// synopsys translate_off
defparam \portA~27 .lut_mask = 16'hCCF0;
defparam \portA~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N0
cycloneive_lcell_comb \portA~28 (
// Equation(s):
// \portA~28_combout  = (fuifforward_A_01 & (!\lui_M~q  & (porto_M_14))) # (!fuifforward_A_01 & (((rdata1_EX[14]))))

	.dataa(\lui_M~q ),
	.datab(porto_M_14),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(rdata1_EX[14]),
	.cin(gnd),
	.combout(\portA~28_combout ),
	.cout());
// synopsys translate_off
defparam \portA~28 .lut_mask = 16'h4F40;
defparam \portA~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N14
cycloneive_lcell_comb \portA~29 (
// Equation(s):
// \portA~29_combout  = (fuifforward_A_11 & (\wdat_WB[14]~37_combout )) # (!fuifforward_A_11 & ((\portA~28_combout )))

	.dataa(\wdat_WB[14]~37_combout ),
	.datab(\portA~28_combout ),
	.datac(gnd),
	.datad(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.cin(gnd),
	.combout(\portA~29_combout ),
	.cout());
// synopsys translate_off
defparam \portA~29 .lut_mask = 16'hAACC;
defparam \portA~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N14
cycloneive_lcell_comb \portA~30 (
// Equation(s):
// \portA~30_combout  = (fuifforward_A_01 & (porto_M_13 & (!\lui_M~q ))) # (!fuifforward_A_01 & (((rdata1_EX[13]))))

	.dataa(porto_M_13),
	.datab(\lui_M~q ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(rdata1_EX[13]),
	.cin(gnd),
	.combout(\portA~30_combout ),
	.cout());
// synopsys translate_off
defparam \portA~30 .lut_mask = 16'h2F20;
defparam \portA~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N20
cycloneive_lcell_comb \portA~31 (
// Equation(s):
// \portA~31_combout  = (fuifforward_A_11 & (\wdat_WB[13]~39_combout )) # (!fuifforward_A_11 & ((\portA~30_combout )))

	.dataa(\wdat_WB[13]~39_combout ),
	.datab(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datac(\portA~30_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\portA~31_combout ),
	.cout());
// synopsys translate_off
defparam \portA~31 .lut_mask = 16'hB8B8;
defparam \portA~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N0
cycloneive_lcell_comb \portA~32 (
// Equation(s):
// \portA~32_combout  = (fuifforward_A_01 & (((porto_M_12 & !\lui_M~q )))) # (!fuifforward_A_01 & (rdata1_EX[12]))

	.dataa(rdata1_EX[12]),
	.datab(porto_M_12),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(\lui_M~q ),
	.cin(gnd),
	.combout(\portA~32_combout ),
	.cout());
// synopsys translate_off
defparam \portA~32 .lut_mask = 16'h0ACA;
defparam \portA~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N2
cycloneive_lcell_comb \portA~33 (
// Equation(s):
// \portA~33_combout  = (fuifforward_A_11 & (\wdat_WB[12]~41_combout )) # (!fuifforward_A_11 & ((\portA~32_combout )))

	.dataa(gnd),
	.datab(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datac(\wdat_WB[12]~41_combout ),
	.datad(\portA~32_combout ),
	.cin(gnd),
	.combout(\portA~33_combout ),
	.cout());
// synopsys translate_off
defparam \portA~33 .lut_mask = 16'hF3C0;
defparam \portA~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N28
cycloneive_lcell_comb \portA~34 (
// Equation(s):
// \portA~34_combout  = (fuifforward_A_01 & (((porto_M_11 & !\lui_M~q )))) # (!fuifforward_A_01 & (rdata1_EX[11]))

	.dataa(rdata1_EX[11]),
	.datab(porto_M_11),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(\lui_M~q ),
	.cin(gnd),
	.combout(\portA~34_combout ),
	.cout());
// synopsys translate_off
defparam \portA~34 .lut_mask = 16'h0ACA;
defparam \portA~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N10
cycloneive_lcell_comb \portA~35 (
// Equation(s):
// \portA~35_combout  = (fuifforward_A_11 & (\wdat_WB[11]~47_combout )) # (!fuifforward_A_11 & ((\portA~34_combout )))

	.dataa(\wdat_WB[11]~47_combout ),
	.datab(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datac(gnd),
	.datad(\portA~34_combout ),
	.cin(gnd),
	.combout(\portA~35_combout ),
	.cout());
// synopsys translate_off
defparam \portA~35 .lut_mask = 16'hBB88;
defparam \portA~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N20
cycloneive_lcell_comb \portA~36 (
// Equation(s):
// \portA~36_combout  = (fuifforward_A_11 & (\wdat_WB[10]~49_combout )) # (!fuifforward_A_11 & ((\portA~71_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[10]~49_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~71_combout ),
	.cin(gnd),
	.combout(\portA~36_combout ),
	.cout());
// synopsys translate_off
defparam \portA~36 .lut_mask = 16'hCFC0;
defparam \portA~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N26
cycloneive_lcell_comb \portA~37 (
// Equation(s):
// \portA~37_combout  = (fuifforward_A_11 & (\wdat_WB[9]~43_combout )) # (!fuifforward_A_11 & ((\portA~72_combout )))

	.dataa(gnd),
	.datab(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datac(\wdat_WB[9]~43_combout ),
	.datad(\portA~72_combout ),
	.cin(gnd),
	.combout(\portA~37_combout ),
	.cout());
// synopsys translate_off
defparam \portA~37 .lut_mask = 16'hF3C0;
defparam \portA~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N18
cycloneive_lcell_comb \portA~38 (
// Equation(s):
// \portA~38_combout  = (fuifforward_A_01 & ((\sw_forwarding_output~0_combout ))) # (!fuifforward_A_01 & (rdata1_EX[31]))

	.dataa(rdata1_EX[31]),
	.datab(gnd),
	.datac(\sw_forwarding_output~0_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~38_combout ),
	.cout());
// synopsys translate_off
defparam \portA~38 .lut_mask = 16'hF0AA;
defparam \portA~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N24
cycloneive_lcell_comb \portA~39 (
// Equation(s):
// \portA~39_combout  = (fuifforward_A_11 & ((\wdat_WB[31]~3_combout ))) # (!fuifforward_A_11 & (\portA~38_combout ))

	.dataa(gnd),
	.datab(\portA~38_combout ),
	.datac(\wdat_WB[31]~3_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.cin(gnd),
	.combout(\portA~39_combout ),
	.cout());
// synopsys translate_off
defparam \portA~39 .lut_mask = 16'hF0CC;
defparam \portA~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N20
cycloneive_lcell_comb \portA~40 (
// Equation(s):
// \portA~40_combout  = (fuifforward_A_01 & ((\sw_forwarding_output~2_combout ))) # (!fuifforward_A_01 & (rdata1_EX[29]))

	.dataa(rdata1_EX[29]),
	.datab(\sw_forwarding_output~2_combout ),
	.datac(gnd),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~40_combout ),
	.cout());
// synopsys translate_off
defparam \portA~40 .lut_mask = 16'hCCAA;
defparam \portA~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N30
cycloneive_lcell_comb \portA~41 (
// Equation(s):
// \portA~41_combout  = (fuifforward_A_11 & (\wdat_WB[29]~7_combout )) # (!fuifforward_A_11 & ((\portA~40_combout )))

	.dataa(gnd),
	.datab(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datac(\wdat_WB[29]~7_combout ),
	.datad(\portA~40_combout ),
	.cin(gnd),
	.combout(\portA~41_combout ),
	.cout());
// synopsys translate_off
defparam \portA~41 .lut_mask = 16'hF3C0;
defparam \portA~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N26
cycloneive_lcell_comb \portA~42 (
// Equation(s):
// \portA~42_combout  = (fuifforward_A_01 & (\sw_forwarding_output~1_combout )) # (!fuifforward_A_01 & ((rdata1_EX[30])))

	.dataa(gnd),
	.datab(\sw_forwarding_output~1_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(rdata1_EX[30]),
	.cin(gnd),
	.combout(\portA~42_combout ),
	.cout());
// synopsys translate_off
defparam \portA~42 .lut_mask = 16'hCFC0;
defparam \portA~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N24
cycloneive_lcell_comb \portA~43 (
// Equation(s):
// \portA~43_combout  = (fuifforward_A_11 & (\wdat_WB[30]~5_combout )) # (!fuifforward_A_11 & ((\portA~42_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[30]~5_combout ),
	.datac(\portA~42_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.cin(gnd),
	.combout(\portA~43_combout ),
	.cout());
// synopsys translate_off
defparam \portA~43 .lut_mask = 16'hCCF0;
defparam \portA~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N10
cycloneive_lcell_comb \portA~44 (
// Equation(s):
// \portA~44_combout  = (fuifforward_A_01 & ((\sw_forwarding_output~3_combout ))) # (!fuifforward_A_01 & (rdata1_EX[28]))

	.dataa(rdata1_EX[28]),
	.datab(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datac(gnd),
	.datad(\sw_forwarding_output~3_combout ),
	.cin(gnd),
	.combout(\portA~44_combout ),
	.cout());
// synopsys translate_off
defparam \portA~44 .lut_mask = 16'hEE22;
defparam \portA~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N22
cycloneive_lcell_comb \portA~45 (
// Equation(s):
// \portA~45_combout  = (fuifforward_A_11 & ((\wdat_WB[28]~9_combout ))) # (!fuifforward_A_11 & (\portA~44_combout ))

	.dataa(\portA~44_combout ),
	.datab(\wdat_WB[28]~9_combout ),
	.datac(gnd),
	.datad(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.cin(gnd),
	.combout(\portA~45_combout ),
	.cout());
// synopsys translate_off
defparam \portA~45 .lut_mask = 16'hCCAA;
defparam \portA~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N16
cycloneive_lcell_comb \portA~46 (
// Equation(s):
// \portA~46_combout  = (fuifforward_A_01 & ((\sw_forwarding_output~4_combout ))) # (!fuifforward_A_01 & (rdata1_EX[27]))

	.dataa(rdata1_EX[27]),
	.datab(\sw_forwarding_output~4_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\portA~46_combout ),
	.cout());
// synopsys translate_off
defparam \portA~46 .lut_mask = 16'hCACA;
defparam \portA~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N22
cycloneive_lcell_comb \portA~47 (
// Equation(s):
// \portA~47_combout  = (fuifforward_A_11 & (\wdat_WB[27]~11_combout )) # (!fuifforward_A_11 & ((\portA~46_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[27]~11_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~46_combout ),
	.cin(gnd),
	.combout(\portA~47_combout ),
	.cout());
// synopsys translate_off
defparam \portA~47 .lut_mask = 16'hCFC0;
defparam \portA~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N18
cycloneive_lcell_comb \portA~48 (
// Equation(s):
// \portA~48_combout  = (fuifforward_A_01 & (\sw_forwarding_output~5_combout )) # (!fuifforward_A_01 & ((rdata1_EX[26])))

	.dataa(gnd),
	.datab(\sw_forwarding_output~5_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(rdata1_EX[26]),
	.cin(gnd),
	.combout(\portA~48_combout ),
	.cout());
// synopsys translate_off
defparam \portA~48 .lut_mask = 16'hCFC0;
defparam \portA~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N12
cycloneive_lcell_comb \portA~49 (
// Equation(s):
// \portA~49_combout  = (fuifforward_A_11 & (\wdat_WB[26]~13_combout )) # (!fuifforward_A_11 & ((\portA~48_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[26]~13_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~48_combout ),
	.cin(gnd),
	.combout(\portA~49_combout ),
	.cout());
// synopsys translate_off
defparam \portA~49 .lut_mask = 16'hCFC0;
defparam \portA~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N22
cycloneive_lcell_comb \portA~50 (
// Equation(s):
// \portA~50_combout  = (fuifforward_A_01 & (\sw_forwarding_output~6_combout )) # (!fuifforward_A_01 & ((rdata1_EX[25])))

	.dataa(\sw_forwarding_output~6_combout ),
	.datab(rdata1_EX[25]),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\portA~50_combout ),
	.cout());
// synopsys translate_off
defparam \portA~50 .lut_mask = 16'hACAC;
defparam \portA~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N0
cycloneive_lcell_comb \portA~51 (
// Equation(s):
// \portA~51_combout  = (fuifforward_A_11 & (\wdat_WB[25]~15_combout )) # (!fuifforward_A_11 & ((\portA~50_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[25]~15_combout ),
	.datac(\portA~50_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.cin(gnd),
	.combout(\portA~51_combout ),
	.cout());
// synopsys translate_off
defparam \portA~51 .lut_mask = 16'hCCF0;
defparam \portA~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N22
cycloneive_lcell_comb \portA~52 (
// Equation(s):
// \portA~52_combout  = (fuifforward_A_01 & (\sw_forwarding_output~7_combout )) # (!fuifforward_A_01 & ((rdata1_EX[24])))

	.dataa(gnd),
	.datab(\sw_forwarding_output~7_combout ),
	.datac(rdata1_EX[24]),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~52_combout ),
	.cout());
// synopsys translate_off
defparam \portA~52 .lut_mask = 16'hCCF0;
defparam \portA~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N0
cycloneive_lcell_comb \portA~53 (
// Equation(s):
// \portA~53_combout  = (fuifforward_A_11 & ((\wdat_WB[24]~17_combout ))) # (!fuifforward_A_11 & (\portA~52_combout ))

	.dataa(gnd),
	.datab(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datac(\portA~52_combout ),
	.datad(\wdat_WB[24]~17_combout ),
	.cin(gnd),
	.combout(\portA~53_combout ),
	.cout());
// synopsys translate_off
defparam \portA~53 .lut_mask = 16'hFC30;
defparam \portA~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N18
cycloneive_lcell_comb \portA~54 (
// Equation(s):
// \portA~54_combout  = (fuifforward_A_01 & (\sw_forwarding_output~8_combout )) # (!fuifforward_A_01 & ((rdata1_EX[23])))

	.dataa(\sw_forwarding_output~8_combout ),
	.datab(rdata1_EX[23]),
	.datac(gnd),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~54_combout ),
	.cout());
// synopsys translate_off
defparam \portA~54 .lut_mask = 16'hAACC;
defparam \portA~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N20
cycloneive_lcell_comb \portA~55 (
// Equation(s):
// \portA~55_combout  = (fuifforward_A_11 & (\wdat_WB[23]~19_combout )) # (!fuifforward_A_11 & ((\portA~54_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[23]~19_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~54_combout ),
	.cin(gnd),
	.combout(\portA~55_combout ),
	.cout());
// synopsys translate_off
defparam \portA~55 .lut_mask = 16'hCFC0;
defparam \portA~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N4
cycloneive_lcell_comb \portA~56 (
// Equation(s):
// \portA~56_combout  = (fuifforward_A_01 & (\sw_forwarding_output~9_combout )) # (!fuifforward_A_01 & ((rdata1_EX[22])))

	.dataa(\sw_forwarding_output~9_combout ),
	.datab(gnd),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(rdata1_EX[22]),
	.cin(gnd),
	.combout(\portA~56_combout ),
	.cout());
// synopsys translate_off
defparam \portA~56 .lut_mask = 16'hAFA0;
defparam \portA~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N8
cycloneive_lcell_comb \portA~57 (
// Equation(s):
// \portA~57_combout  = (fuifforward_A_11 & (\wdat_WB[22]~21_combout )) # (!fuifforward_A_11 & ((\portA~56_combout )))

	.dataa(gnd),
	.datab(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datac(\wdat_WB[22]~21_combout ),
	.datad(\portA~56_combout ),
	.cin(gnd),
	.combout(\portA~57_combout ),
	.cout());
// synopsys translate_off
defparam \portA~57 .lut_mask = 16'hF3C0;
defparam \portA~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N2
cycloneive_lcell_comb \portA~58 (
// Equation(s):
// \portA~58_combout  = (fuifforward_A_01 & ((\sw_forwarding_output~10_combout ))) # (!fuifforward_A_01 & (rdata1_EX[21]))

	.dataa(rdata1_EX[21]),
	.datab(\sw_forwarding_output~10_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\portA~58_combout ),
	.cout());
// synopsys translate_off
defparam \portA~58 .lut_mask = 16'hCACA;
defparam \portA~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N12
cycloneive_lcell_comb \portA~59 (
// Equation(s):
// \portA~59_combout  = (fuifforward_A_11 & (\wdat_WB[21]~23_combout )) # (!fuifforward_A_11 & ((\portA~58_combout )))

	.dataa(gnd),
	.datab(\wdat_WB[21]~23_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~58_combout ),
	.cin(gnd),
	.combout(\portA~59_combout ),
	.cout());
// synopsys translate_off
defparam \portA~59 .lut_mask = 16'hCFC0;
defparam \portA~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N0
cycloneive_lcell_comb \portA~60 (
// Equation(s):
// \portA~60_combout  = (fuifforward_A_01 & (\sw_forwarding_output~11_combout )) # (!fuifforward_A_01 & ((rdata1_EX[20])))

	.dataa(gnd),
	.datab(\sw_forwarding_output~11_combout ),
	.datac(rdata1_EX[20]),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~60_combout ),
	.cout());
// synopsys translate_off
defparam \portA~60 .lut_mask = 16'hCCF0;
defparam \portA~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N30
cycloneive_lcell_comb \portA~61 (
// Equation(s):
// \portA~61_combout  = (fuifforward_A_11 & (\wdat_WB[20]~25_combout )) # (!fuifforward_A_11 & ((\portA~60_combout )))

	.dataa(\wdat_WB[20]~25_combout ),
	.datab(gnd),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~60_combout ),
	.cin(gnd),
	.combout(\portA~61_combout ),
	.cout());
// synopsys translate_off
defparam \portA~61 .lut_mask = 16'hAFA0;
defparam \portA~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N20
cycloneive_lcell_comb \portA~62 (
// Equation(s):
// \portA~62_combout  = (fuifforward_A_01 & (\sw_forwarding_output~12_combout )) # (!fuifforward_A_01 & ((rdata1_EX[19])))

	.dataa(gnd),
	.datab(\sw_forwarding_output~12_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(rdata1_EX[19]),
	.cin(gnd),
	.combout(\portA~62_combout ),
	.cout());
// synopsys translate_off
defparam \portA~62 .lut_mask = 16'hCFC0;
defparam \portA~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N30
cycloneive_lcell_comb \portA~63 (
// Equation(s):
// \portA~63_combout  = (fuifforward_A_11 & ((\wdat_WB[19]~27_combout ))) # (!fuifforward_A_11 & (\portA~62_combout ))

	.dataa(gnd),
	.datab(\portA~62_combout ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\wdat_WB[19]~27_combout ),
	.cin(gnd),
	.combout(\portA~63_combout ),
	.cout());
// synopsys translate_off
defparam \portA~63 .lut_mask = 16'hFC0C;
defparam \portA~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N12
cycloneive_lcell_comb \portA~64 (
// Equation(s):
// \portA~64_combout  = (fuifforward_A_01 & ((\sw_forwarding_output~13_combout ))) # (!fuifforward_A_01 & (rdata1_EX[18]))

	.dataa(rdata1_EX[18]),
	.datab(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datac(gnd),
	.datad(\sw_forwarding_output~13_combout ),
	.cin(gnd),
	.combout(\portA~64_combout ),
	.cout());
// synopsys translate_off
defparam \portA~64 .lut_mask = 16'hEE22;
defparam \portA~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N14
cycloneive_lcell_comb \portA~65 (
// Equation(s):
// \portA~65_combout  = (fuifforward_A_11 & ((\wdat_WB[18]~29_combout ))) # (!fuifforward_A_11 & (\portA~64_combout ))

	.dataa(\portA~64_combout ),
	.datab(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datac(gnd),
	.datad(\wdat_WB[18]~29_combout ),
	.cin(gnd),
	.combout(\portA~65_combout ),
	.cout());
// synopsys translate_off
defparam \portA~65 .lut_mask = 16'hEE22;
defparam \portA~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N24
cycloneive_lcell_comb \portA~66 (
// Equation(s):
// \portA~66_combout  = (fuifforward_A_01 & ((\sw_forwarding_output~14_combout ))) # (!fuifforward_A_01 & (rdata1_EX[17]))

	.dataa(gnd),
	.datab(rdata1_EX[17]),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(\sw_forwarding_output~14_combout ),
	.cin(gnd),
	.combout(\portA~66_combout ),
	.cout());
// synopsys translate_off
defparam \portA~66 .lut_mask = 16'hFC0C;
defparam \portA~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N10
cycloneive_lcell_comb \portA~67 (
// Equation(s):
// \portA~67_combout  = (fuifforward_A_11 & (\wdat_WB[17]~31_combout )) # (!fuifforward_A_11 & ((\portA~66_combout )))

	.dataa(\wdat_WB[17]~31_combout ),
	.datab(gnd),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\portA~66_combout ),
	.cin(gnd),
	.combout(\portA~67_combout ),
	.cout());
// synopsys translate_off
defparam \portA~67 .lut_mask = 16'hAFA0;
defparam \portA~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N17
dffeas \btbframes.frameblocks[2].jump_add[1] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N23
dffeas \btbframes.frameblocks[1].jump_add[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N29
dffeas \btbframes.frameblocks[0].jump_add[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N28
cycloneive_lcell_comb \pc_next[1]~0 (
// Equation(s):
// \pc_next[1]~0_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].jump_add [1])) # (!pc_out_2 & ((\btbframes.frameblocks[0].jump_add [1])))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[1].jump_add [1]),
	.datac(\btbframes.frameblocks[0].jump_add [1]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[1]~0 .lut_mask = 16'hEE50;
defparam \pc_next[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N31
dffeas \btbframes.frameblocks[3].jump_add[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N30
cycloneive_lcell_comb \pc_next[1]~1 (
// Equation(s):
// \pc_next[1]~1_combout  = (\pc_next[1]~0_combout  & (((\btbframes.frameblocks[3].jump_add [1])) # (!pc_out_3))) # (!\pc_next[1]~0_combout  & (pc_out_3 & ((\btbframes.frameblocks[2].jump_add [1]))))

	.dataa(\pc_next[1]~0_combout ),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[3].jump_add [1]),
	.datad(\btbframes.frameblocks[2].jump_add [1]),
	.cin(gnd),
	.combout(\pc_next[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[1]~1 .lut_mask = 16'hE6A2;
defparam \pc_next[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N4
cycloneive_lcell_comb \pc_next[1]~2 (
// Equation(s):
// \pc_next[1]~2_combout  = (\jr_M~q  & ((rdata1_M[1]))) # (!\jr_M~q  & (pc_plus_4_M[1]))

	.dataa(pc_plus_4_M[1]),
	.datab(gnd),
	.datac(rdata1_M[1]),
	.datad(\jr_M~q ),
	.cin(gnd),
	.combout(\pc_next[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[1]~2 .lut_mask = 16'hF0AA;
defparam \pc_next[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N9
dffeas \btbframes.frameblocks[2].tag[1] (
	.clk(CLK),
	.d(\Add2~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N25
dffeas \btbframes.frameblocks[1].tag[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N1
dffeas \btbframes.frameblocks[0].tag[1] (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].tag[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N31
dffeas \btbframes.frameblocks[3].tag[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N1
dffeas \btbframes.frameblocks[1].tag[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N1
dffeas \btbframes.frameblocks[2].tag[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N19
dffeas \btbframes.frameblocks[0].tag[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N7
dffeas \btbframes.frameblocks[3].tag[0] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N17
dffeas \btbframes.frameblocks[2].tag[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [3]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[3] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N13
dffeas \btbframes.frameblocks[1].tag[3] (
	.clk(CLK),
	.d(\Add2~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [3]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[3] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N3
dffeas \btbframes.frameblocks[0].tag[3] (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].tag[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [3]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[3] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N5
dffeas \btbframes.frameblocks[3].tag[3] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [3]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[3] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N11
dffeas \btbframes.frameblocks[1].tag[2] (
	.clk(CLK),
	.d(\Add2~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [2]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[2] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N23
dffeas \btbframes.frameblocks[2].tag[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [2]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[2] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y40_N29
dffeas \btbframes.frameblocks[0].tag[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [2]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[2] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N21
dffeas \btbframes.frameblocks[3].tag[2] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [2]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[2] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N19
dffeas \btbframes.frameblocks[2].tag[5] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].tag[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [5]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[5] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N17
dffeas \btbframes.frameblocks[1].tag[5] (
	.clk(CLK),
	.d(\Add2~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [5]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[5] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N1
dffeas \btbframes.frameblocks[0].tag[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [5]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[5] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N3
dffeas \btbframes.frameblocks[3].tag[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [5]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[5] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N15
dffeas \btbframes.frameblocks[1].tag[4] (
	.clk(CLK),
	.d(\Add2~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [4]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[4] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N7
dffeas \btbframes.frameblocks[2].tag[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [4]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[4] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N5
dffeas \btbframes.frameblocks[0].tag[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [4]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[4] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N25
dffeas \btbframes.frameblocks[3].tag[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [4]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[4] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N21
dffeas \btbframes.frameblocks[2].tag[7] (
	.clk(CLK),
	.d(\Add2~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [7]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[7] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N1
dffeas \btbframes.frameblocks[1].tag[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [7]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[7] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N7
dffeas \btbframes.frameblocks[0].tag[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [7]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[7] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N29
dffeas \btbframes.frameblocks[3].tag[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [7]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[7] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N15
dffeas \btbframes.frameblocks[1].tag[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [6]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[6] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N19
dffeas \btbframes.frameblocks[2].tag[6] (
	.clk(CLK),
	.d(\Add2~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [6]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[6] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N31
dffeas \btbframes.frameblocks[0].tag[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [6]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[6] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N1
dffeas \btbframes.frameblocks[3].tag[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [6]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[6] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N11
dffeas \btbframes.frameblocks[2].tag[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [9]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[9] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N17
dffeas \btbframes.frameblocks[1].tag[9] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].tag[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [9]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[9] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N25
dffeas \btbframes.frameblocks[0].tag[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [9]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[9] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N11
dffeas \btbframes.frameblocks[3].tag[9] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [9]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[9] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N27
dffeas \btbframes.frameblocks[1].tag[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [8]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[8] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N21
dffeas \btbframes.frameblocks[2].tag[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [8]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[8] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N11
dffeas \btbframes.frameblocks[0].tag[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [8]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[8] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N17
dffeas \btbframes.frameblocks[3].tag[8] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [8]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[8] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N29
dffeas \btbframes.frameblocks[2].tag[11] (
	.clk(CLK),
	.d(\Add2~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [11]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[11] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N7
dffeas \btbframes.frameblocks[1].tag[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [11]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[11] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N29
dffeas \btbframes.frameblocks[0].tag[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [11]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[11] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N17
dffeas \btbframes.frameblocks[3].tag[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [11]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[11] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N13
dffeas \btbframes.frameblocks[1].tag[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [10]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[10] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N15
dffeas \btbframes.frameblocks[2].tag[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [10]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[10] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N13
dffeas \btbframes.frameblocks[0].tag[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [10]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[10] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N3
dffeas \btbframes.frameblocks[3].tag[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [10]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[10] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N1
dffeas \btbframes.frameblocks[2].tag[13] (
	.clk(CLK),
	.d(\Add2~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [13]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[13] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N15
dffeas \btbframes.frameblocks[1].tag[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [13]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[13] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N27
dffeas \btbframes.frameblocks[0].tag[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [13]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[13] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N21
dffeas \btbframes.frameblocks[3].tag[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [13]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[13] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N7
dffeas \btbframes.frameblocks[1].tag[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [12]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[12] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N23
dffeas \btbframes.frameblocks[2].tag[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [12]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[12] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N5
dffeas \btbframes.frameblocks[0].tag[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [12]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[12] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N25
dffeas \btbframes.frameblocks[3].tag[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [12]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[12] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N15
dffeas \btbframes.frameblocks[2].tag[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~34_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [15]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[15] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N3
dffeas \btbframes.frameblocks[1].tag[15] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].tag[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [15]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[15] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N5
dffeas \btbframes.frameblocks[0].tag[15] (
	.clk(CLK),
	.d(\Add2~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [15]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[15] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N27
dffeas \btbframes.frameblocks[3].tag[15] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [15]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[15] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N13
dffeas \btbframes.frameblocks[1].tag[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [14]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[14] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N27
dffeas \btbframes.frameblocks[2].tag[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [14]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[14] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N25
dffeas \btbframes.frameblocks[0].tag[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [14]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[14] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y39_N23
dffeas \btbframes.frameblocks[3].tag[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [14]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[14] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N9
dffeas \btbframes.frameblocks[2].tag[17] (
	.clk(CLK),
	.d(\Add2~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [17]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[17] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N1
dffeas \btbframes.frameblocks[1].tag[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~38_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [17]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[17] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N3
dffeas \btbframes.frameblocks[0].tag[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~38_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [17]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[17] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N23
dffeas \btbframes.frameblocks[3].tag[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~38_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [17]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[17] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N9
dffeas \btbframes.frameblocks[1].tag[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~36_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [16]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[16] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y41_N17
dffeas \btbframes.frameblocks[2].tag[16] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].tag[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [16]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[16] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N7
dffeas \btbframes.frameblocks[0].tag[16] (
	.clk(CLK),
	.d(\Add2~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [16]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[16] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N5
dffeas \btbframes.frameblocks[3].tag[16] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [16]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[16] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N5
dffeas \btbframes.frameblocks[2].tag[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [19]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[19] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N25
dffeas \btbframes.frameblocks[1].tag[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [19]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[19] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N21
dffeas \btbframes.frameblocks[0].tag[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [19]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[19] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N31
dffeas \btbframes.frameblocks[3].tag[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [19]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[19] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N1
dffeas \btbframes.frameblocks[1].tag[18] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].tag[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [18]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[18] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N13
dffeas \btbframes.frameblocks[2].tag[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~40_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [18]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[18] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N11
dffeas \btbframes.frameblocks[0].tag[18] (
	.clk(CLK),
	.d(\Add2~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [18]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[18] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N29
dffeas \btbframes.frameblocks[3].tag[18] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [18]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[18] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y39_N7
dffeas \btbframes.frameblocks[2].tag[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [21]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[21] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N31
dffeas \btbframes.frameblocks[1].tag[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [21]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[21] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N3
dffeas \btbframes.frameblocks[0].tag[21] (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].tag[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [21]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[21] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N17
dffeas \btbframes.frameblocks[3].tag[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [21]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[21] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N27
dffeas \btbframes.frameblocks[1].tag[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~44_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [20]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[20] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N31
dffeas \btbframes.frameblocks[2].tag[20] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].tag[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [20]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[20] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y40_N7
dffeas \btbframes.frameblocks[0].tag[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~44_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [20]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[20] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N21
dffeas \btbframes.frameblocks[3].tag[20] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [20]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[20] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N21
dffeas \btbframes.frameblocks[2].tag[23] (
	.clk(CLK),
	.d(\Add2~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [23]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[23] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N23
dffeas \btbframes.frameblocks[1].tag[23] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].tag[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [23]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[23] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N13
dffeas \btbframes.frameblocks[0].tag[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~50_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [23]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[23] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N15
dffeas \btbframes.frameblocks[3].tag[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~50_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [23]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[23] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N1
dffeas \btbframes.frameblocks[1].tag[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~48_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [22]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[22] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N3
dffeas \btbframes.frameblocks[2].tag[22] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].tag[22]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [22]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[22] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N19
dffeas \btbframes.frameblocks[0].tag[22] (
	.clk(CLK),
	.d(\Add2~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [22]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[22] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N27
dffeas \btbframes.frameblocks[3].tag[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~48_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [22]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[22] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N25
dffeas \btbframes.frameblocks[2].tag[25] (
	.clk(CLK),
	.d(\Add2~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [25]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[25] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N25
dffeas \btbframes.frameblocks[1].tag[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [25]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[25] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N13
dffeas \btbframes.frameblocks[0].tag[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [25]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[25] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N23
dffeas \btbframes.frameblocks[3].tag[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [25]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[25] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N9
dffeas \btbframes.frameblocks[1].tag[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [24]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[24] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N9
dffeas \btbframes.frameblocks[2].tag[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [24]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[24] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N31
dffeas \btbframes.frameblocks[0].tag[24] (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].tag[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [24]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[24] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N19
dffeas \btbframes.frameblocks[3].tag[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [24]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[24] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N11
dffeas \btbframes.frameblocks[2].tag[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [27]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[27] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N23
dffeas \btbframes.frameblocks[1].tag[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [27]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[27] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N17
dffeas \btbframes.frameblocks[0].tag[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [27]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[27] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N29
dffeas \btbframes.frameblocks[3].tag[27] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[27]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [27]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[27] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N25
dffeas \btbframes.frameblocks[1].tag[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~56_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].tag [26]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[26] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].tag[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N1
dffeas \btbframes.frameblocks[2].tag[26] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].tag[26]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].tag [26]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[26] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].tag[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N13
dffeas \btbframes.frameblocks[0].tag[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Add2~56_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].tag [26]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[26] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].tag[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N27
dffeas \btbframes.frameblocks[3].tag[26] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].tag[26]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].tag [26]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[26] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].tag[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N3
dffeas \btbframes.frameblocks[2].valid (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].valid~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].valid~q ),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].valid .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].valid .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N21
dffeas \btbframes.frameblocks[1].valid (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].valid~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].valid~q ),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].valid .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].valid .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N27
dffeas \btbframes.frameblocks[0].valid (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].valid~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].valid~q ),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].valid .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].valid .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y40_N15
dffeas \btbframes.frameblocks[3].valid (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].valid~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].valid~q ),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].valid .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].valid .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N5
dffeas \btbframes.frameblocks[1].curr_state[1] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].curr_state[1]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].curr_state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].curr_state[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].curr_state[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N7
dffeas \btbframes.frameblocks[2].curr_state[1] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].curr_state[1]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].curr_state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].curr_state[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].curr_state[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N29
dffeas \btbframes.frameblocks[0].curr_state[1] (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].curr_state[1]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].curr_state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].curr_state[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].curr_state[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N23
dffeas \btbframes.frameblocks[3].curr_state[1] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].curr_state[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].curr_state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].curr_state[1] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].curr_state[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N30
cycloneive_lcell_comb \pc_next~3 (
// Equation(s):
// \pc_next~3_combout  = (\branch_or_jump~1_combout  & predicted)

	.dataa(gnd),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\BTB|predicted~18_combout ),
	.cin(gnd),
	.combout(\pc_next~3_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next~3 .lut_mask = 16'hF000;
defparam \pc_next~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N28
cycloneive_lcell_comb \pc_next[1]~4 (
// Equation(s):
// \pc_next[1]~4_combout  = (\pc_next~3_combout  & (((\pc_next[1]~1_combout )))) # (!\pc_next~3_combout  & (\pc_next[1]~2_combout  & (\branch_or_jump~0_combout )))

	.dataa(\pc_next[1]~2_combout ),
	.datab(\branch_or_jump~0_combout ),
	.datac(\pc_next[1]~1_combout ),
	.datad(\pc_next~3_combout ),
	.cin(gnd),
	.combout(\pc_next[1]~4_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[1]~4 .lut_mask = 16'hF088;
defparam \pc_next[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N22
cycloneive_lcell_comb \portB~108 (
// Equation(s):
// \portB~108_combout  = (\portB~78_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(\Equal3~2_combout ),
	.datab(\ShiftOp_EX~q ),
	.datac(gnd),
	.datad(\portB~78_combout ),
	.cin(gnd),
	.combout(\portB~108_combout ),
	.cout());
// synopsys translate_off
defparam \portB~108 .lut_mask = 16'hBB00;
defparam \portB~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N28
cycloneive_lcell_comb \portB~109 (
// Equation(s):
// \portB~109_combout  = (\portB~80_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(gnd),
	.datab(\ShiftOp_EX~q ),
	.datac(\Equal3~2_combout ),
	.datad(\portB~80_combout ),
	.cin(gnd),
	.combout(\portB~109_combout ),
	.cout());
// synopsys translate_off
defparam \portB~109 .lut_mask = 16'hF300;
defparam \portB~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N13
dffeas \btbframes.frameblocks[1].jump_add[0] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N1
dffeas \btbframes.frameblocks[2].jump_add[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[0]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N23
dffeas \btbframes.frameblocks[0].jump_add[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[0]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N22
cycloneive_lcell_comb \pc_next[0]~5 (
// Equation(s):
// \pc_next[0]~5_combout  = (pc_out_2 & (pc_out_3)) # (!pc_out_2 & ((pc_out_3 & ((\btbframes.frameblocks[2].jump_add [0]))) # (!pc_out_3 & (\btbframes.frameblocks[0].jump_add [0]))))

	.dataa(pc_out_2),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[0].jump_add [0]),
	.datad(\btbframes.frameblocks[2].jump_add [0]),
	.cin(gnd),
	.combout(\pc_next[0]~5_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[0]~5 .lut_mask = 16'hDC98;
defparam \pc_next[0]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N19
dffeas \btbframes.frameblocks[3].jump_add[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[0]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N18
cycloneive_lcell_comb \pc_next[0]~6 (
// Equation(s):
// \pc_next[0]~6_combout  = (pc_out_2 & ((\pc_next[0]~5_combout  & ((\btbframes.frameblocks[3].jump_add [0]))) # (!\pc_next[0]~5_combout  & (\btbframes.frameblocks[1].jump_add [0])))) # (!pc_out_2 & (((\pc_next[0]~5_combout ))))

	.dataa(\btbframes.frameblocks[1].jump_add [0]),
	.datab(pc_out_2),
	.datac(\btbframes.frameblocks[3].jump_add [0]),
	.datad(\pc_next[0]~5_combout ),
	.cin(gnd),
	.combout(\pc_next[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[0]~6 .lut_mask = 16'hF388;
defparam \pc_next[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N14
cycloneive_lcell_comb \pc_next[0]~7 (
// Equation(s):
// \pc_next[0]~7_combout  = (\jr_M~q  & (rdata1_M[0])) # (!\jr_M~q  & ((pc_plus_4_M[0])))

	.dataa(\jr_M~q ),
	.datab(gnd),
	.datac(rdata1_M[0]),
	.datad(pc_plus_4_M[0]),
	.cin(gnd),
	.combout(\pc_next[0]~7_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[0]~7 .lut_mask = 16'hF5A0;
defparam \pc_next[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N22
cycloneive_lcell_comb \pc_next[0]~8 (
// Equation(s):
// \pc_next[0]~8_combout  = (\pc_next~3_combout  & (((\pc_next[0]~6_combout )))) # (!\pc_next~3_combout  & (\branch_or_jump~0_combout  & ((\pc_next[0]~7_combout ))))

	.dataa(\branch_or_jump~0_combout ),
	.datab(\pc_next[0]~6_combout ),
	.datac(\pc_next[0]~7_combout ),
	.datad(\pc_next~3_combout ),
	.cin(gnd),
	.combout(\pc_next[0]~8_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[0]~8 .lut_mask = 16'hCCA0;
defparam \pc_next[0]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N20
cycloneive_lcell_comb \pc_next[3]~9 (
// Equation(s):
// \pc_next[3]~9_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & (\pc_when_branch[3]~2_combout )) # (!pc_out_101 & ((pc_plus_4_M[3]))))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(\pc_when_branch[3]~2_combout ),
	.datab(\branch_or_jump~2_combout ),
	.datac(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datad(pc_plus_4_M[3]),
	.cin(gnd),
	.combout(\pc_next[3]~9_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[3]~9 .lut_mask = 16'hBCB0;
defparam \pc_next[3]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N2
cycloneive_lcell_comb \pc_next[3]~10 (
// Equation(s):
// \pc_next[3]~10_combout  = (\branch_or_jump~2_combout  & (((\pc_next[3]~9_combout )))) # (!\branch_or_jump~2_combout  & ((\pc_next[3]~9_combout  & (imm_M[1])) # (!\pc_next[3]~9_combout  & ((rdata1_M[3])))))

	.dataa(imm_M[1]),
	.datab(\branch_or_jump~2_combout ),
	.datac(rdata1_M[3]),
	.datad(\pc_next[3]~9_combout ),
	.cin(gnd),
	.combout(\pc_next[3]~10_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[3]~10 .lut_mask = 16'hEE30;
defparam \pc_next[3]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N9
dffeas \btbframes.frameblocks[1].jump_add[3] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [3]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[3] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N25
dffeas \btbframes.frameblocks[2].jump_add[3] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [3]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[3] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N7
dffeas \btbframes.frameblocks[0].jump_add[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[3]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [3]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[3] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N6
cycloneive_lcell_comb \pc_next[3]~11 (
// Equation(s):
// \pc_next[3]~11_combout  = (pc_out_3 & ((\btbframes.frameblocks[2].jump_add [3]) # ((pc_out_2)))) # (!pc_out_3 & (((\btbframes.frameblocks[0].jump_add [3] & !pc_out_2))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[2].jump_add [3]),
	.datac(\btbframes.frameblocks[0].jump_add [3]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[3]~11_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[3]~11 .lut_mask = 16'hAAD8;
defparam \pc_next[3]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N31
dffeas \btbframes.frameblocks[3].jump_add[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[3]~2_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [3]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[3] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N30
cycloneive_lcell_comb \pc_next[3]~12 (
// Equation(s):
// \pc_next[3]~12_combout  = (\pc_next[3]~11_combout  & (((\btbframes.frameblocks[3].jump_add [3])) # (!pc_out_2))) # (!\pc_next[3]~11_combout  & (pc_out_2 & ((\btbframes.frameblocks[1].jump_add [3]))))

	.dataa(\pc_next[3]~11_combout ),
	.datab(pc_out_2),
	.datac(\btbframes.frameblocks[3].jump_add [3]),
	.datad(\btbframes.frameblocks[1].jump_add [3]),
	.cin(gnd),
	.combout(\pc_next[3]~12_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[3]~12 .lut_mask = 16'hE6A2;
defparam \pc_next[3]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N18
cycloneive_lcell_comb \comb~2 (
// Equation(s):
// \comb~2_combout  = ((!dhit & (always1 & !Decoder11))) # (!\branch_or_jump~1_combout )

	.dataa(dhit),
	.datab(\branch_or_jump~1_combout ),
	.datac(always1),
	.datad(\CONTROL_UNIT|Decoder1~1_combout ),
	.cin(gnd),
	.combout(\comb~2_combout ),
	.cout());
// synopsys translate_off
defparam \comb~2 .lut_mask = 16'h3373;
defparam \comb~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N28
cycloneive_lcell_comb \pc_next[2]~13 (
// Equation(s):
// \pc_next[2]~13_combout  = (\branch_or_jump~2_combout  & (!pc_out_101 & (pc_plus_4_M[2]))) # (!\branch_or_jump~2_combout  & ((pc_out_101) # ((rdata1_M[2]))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datac(pc_plus_4_M[2]),
	.datad(rdata1_M[2]),
	.cin(gnd),
	.combout(\pc_next[2]~13_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[2]~13 .lut_mask = 16'h7564;
defparam \pc_next[2]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N18
cycloneive_lcell_comb \pc_next[2]~14 (
// Equation(s):
// \pc_next[2]~14_combout  = (pc_out_101 & ((\pc_next[2]~13_combout  & (imm_M[0])) # (!\pc_next[2]~13_combout  & ((\pc_when_branch[2]~0_combout ))))) # (!pc_out_101 & (((\pc_next[2]~13_combout ))))

	.dataa(imm_M[0]),
	.datab(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datac(\pc_when_branch[2]~0_combout ),
	.datad(\pc_next[2]~13_combout ),
	.cin(gnd),
	.combout(\pc_next[2]~14_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[2]~14 .lut_mask = 16'hBBC0;
defparam \pc_next[2]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N3
dffeas \btbframes.frameblocks[2].jump_add[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[2]~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [2]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[2] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y41_N25
dffeas \btbframes.frameblocks[1].jump_add[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[2]~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [2]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[2] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N15
dffeas \btbframes.frameblocks[0].jump_add[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[2]~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [2]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[2] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N24
cycloneive_lcell_comb \pc_next[2]~15 (
// Equation(s):
// \pc_next[2]~15_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & ((\btbframes.frameblocks[1].jump_add [2]))) # (!pc_out_2 & (\btbframes.frameblocks[0].jump_add [2]))))

	.dataa(\btbframes.frameblocks[0].jump_add [2]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[1].jump_add [2]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[2]~15_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[2]~15 .lut_mask = 16'hFC22;
defparam \pc_next[2]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y41_N3
dffeas \btbframes.frameblocks[3].jump_add[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[2]~0_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [2]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[2] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N2
cycloneive_lcell_comb \pc_next[2]~16 (
// Equation(s):
// \pc_next[2]~16_combout  = (pc_out_3 & ((\pc_next[2]~15_combout  & ((\btbframes.frameblocks[3].jump_add [2]))) # (!\pc_next[2]~15_combout  & (\btbframes.frameblocks[2].jump_add [2])))) # (!pc_out_3 & (((\pc_next[2]~15_combout ))))

	.dataa(\btbframes.frameblocks[2].jump_add [2]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[3].jump_add [2]),
	.datad(\pc_next[2]~15_combout ),
	.cin(gnd),
	.combout(\pc_next[2]~16_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[2]~16 .lut_mask = 16'hF388;
defparam \pc_next[2]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N18
cycloneive_lcell_comb \pc_next[5]~17 (
// Equation(s):
// \pc_next[5]~17_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_M[5] & (!pc_out_101))) # (!\branch_or_jump~2_combout  & (((pc_out_101) # (rdata1_M[5]))))

	.dataa(pc_plus_4_M[5]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datad(rdata1_M[5]),
	.cin(gnd),
	.combout(\pc_next[5]~17_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[5]~17 .lut_mask = 16'h3B38;
defparam \pc_next[5]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N24
cycloneive_lcell_comb \pc_next[5]~18 (
// Equation(s):
// \pc_next[5]~18_combout  = (\pc_next[5]~17_combout  & (((imm_M[3])) # (!pc_out_101))) # (!\pc_next[5]~17_combout  & (pc_out_101 & ((\pc_when_branch[5]~6_combout ))))

	.dataa(\pc_next[5]~17_combout ),
	.datab(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datac(imm_M[3]),
	.datad(\pc_when_branch[5]~6_combout ),
	.cin(gnd),
	.combout(\pc_next[5]~18_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[5]~18 .lut_mask = 16'hE6A2;
defparam \pc_next[5]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N9
dffeas \btbframes.frameblocks[2].jump_add[5] (
	.clk(CLK),
	.d(\pc_when_branch[5]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [5]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[5] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N9
dffeas \btbframes.frameblocks[1].jump_add[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[5]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [5]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[5] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N1
dffeas \btbframes.frameblocks[0].jump_add[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[5]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [5]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[5] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N0
cycloneive_lcell_comb \pc_next[5]~19 (
// Equation(s):
// \pc_next[5]~19_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].jump_add [5])) # (!pc_out_2 & ((\btbframes.frameblocks[0].jump_add [5])))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[1].jump_add [5]),
	.datac(\btbframes.frameblocks[0].jump_add [5]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[5]~19_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[5]~19 .lut_mask = 16'hEE50;
defparam \pc_next[5]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N27
dffeas \btbframes.frameblocks[3].jump_add[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[5]~6_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [5]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[5] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N26
cycloneive_lcell_comb \pc_next[5]~20 (
// Equation(s):
// \pc_next[5]~20_combout  = (pc_out_3 & ((\pc_next[5]~19_combout  & (\btbframes.frameblocks[3].jump_add [5])) # (!\pc_next[5]~19_combout  & ((\btbframes.frameblocks[2].jump_add [5]))))) # (!pc_out_3 & (\pc_next[5]~19_combout ))

	.dataa(pc_out_3),
	.datab(\pc_next[5]~19_combout ),
	.datac(\btbframes.frameblocks[3].jump_add [5]),
	.datad(\btbframes.frameblocks[2].jump_add [5]),
	.cin(gnd),
	.combout(\pc_next[5]~20_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[5]~20 .lut_mask = 16'hE6C4;
defparam \pc_next[5]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N20
cycloneive_lcell_comb \pc_next[4]~21 (
// Equation(s):
// \pc_next[4]~21_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & ((\pc_when_branch[4]~4_combout ))) # (!pc_out_101 & (pc_plus_4_M[4])))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_M[4]),
	.datac(\pc_when_branch[4]~4_combout ),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[4]~21_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[4]~21 .lut_mask = 16'hF588;
defparam \pc_next[4]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N22
cycloneive_lcell_comb \pc_next[4]~22 (
// Equation(s):
// \pc_next[4]~22_combout  = (\pc_next[4]~21_combout  & ((imm_M[2]) # ((\branch_or_jump~2_combout )))) # (!\pc_next[4]~21_combout  & (((!\branch_or_jump~2_combout  & rdata1_M[4]))))

	.dataa(imm_M[2]),
	.datab(\pc_next[4]~21_combout ),
	.datac(\branch_or_jump~2_combout ),
	.datad(rdata1_M[4]),
	.cin(gnd),
	.combout(\pc_next[4]~22_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[4]~22 .lut_mask = 16'hCBC8;
defparam \pc_next[4]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N29
dffeas \btbframes.frameblocks[1].jump_add[4] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [4]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[4] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N7
dffeas \btbframes.frameblocks[2].jump_add[4] (
	.clk(CLK),
	.d(\pc_when_branch[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [4]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[4] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N29
dffeas \btbframes.frameblocks[0].jump_add[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[4]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [4]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[4] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N28
cycloneive_lcell_comb \pc_next[4]~23 (
// Equation(s):
// \pc_next[4]~23_combout  = (pc_out_2 & (pc_out_3)) # (!pc_out_2 & ((pc_out_3 & ((\btbframes.frameblocks[2].jump_add [4]))) # (!pc_out_3 & (\btbframes.frameblocks[0].jump_add [4]))))

	.dataa(pc_out_2),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[0].jump_add [4]),
	.datad(\btbframes.frameblocks[2].jump_add [4]),
	.cin(gnd),
	.combout(\pc_next[4]~23_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[4]~23 .lut_mask = 16'hDC98;
defparam \pc_next[4]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N11
dffeas \btbframes.frameblocks[3].jump_add[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[4]~4_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [4]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[4] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N10
cycloneive_lcell_comb \pc_next[4]~24 (
// Equation(s):
// \pc_next[4]~24_combout  = (\pc_next[4]~23_combout  & (((\btbframes.frameblocks[3].jump_add [4]) # (!pc_out_2)))) # (!\pc_next[4]~23_combout  & (\btbframes.frameblocks[1].jump_add [4] & ((pc_out_2))))

	.dataa(\pc_next[4]~23_combout ),
	.datab(\btbframes.frameblocks[1].jump_add [4]),
	.datac(\btbframes.frameblocks[3].jump_add [4]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[4]~24_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[4]~24 .lut_mask = 16'hE4AA;
defparam \pc_next[4]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N12
cycloneive_lcell_comb \pc_next[7]~25 (
// Equation(s):
// \pc_next[7]~25_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_M[7] & (!pc_out_101))) # (!\branch_or_jump~2_combout  & (((pc_out_101) # (rdata1_M[7]))))

	.dataa(pc_plus_4_M[7]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datad(rdata1_M[7]),
	.cin(gnd),
	.combout(\pc_next[7]~25_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[7]~25 .lut_mask = 16'h3B38;
defparam \pc_next[7]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N10
cycloneive_lcell_comb \pc_next[7]~26 (
// Equation(s):
// \pc_next[7]~26_combout  = (\pc_next[7]~25_combout  & (((imm_M[5]) # (!pc_out_101)))) # (!\pc_next[7]~25_combout  & (\pc_when_branch[7]~10_combout  & (pc_out_101)))

	.dataa(\pc_next[7]~25_combout ),
	.datab(\pc_when_branch[7]~10_combout ),
	.datac(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datad(imm_M[5]),
	.cin(gnd),
	.combout(\pc_next[7]~26_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[7]~26 .lut_mask = 16'hEA4A;
defparam \pc_next[7]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N9
dffeas \btbframes.frameblocks[2].jump_add[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[7]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [7]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[7] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N11
dffeas \btbframes.frameblocks[1].jump_add[7] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [7]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[7] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N19
dffeas \btbframes.frameblocks[0].jump_add[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[7]~10_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [7]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[7] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N18
cycloneive_lcell_comb \pc_next[7]~27 (
// Equation(s):
// \pc_next[7]~27_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].jump_add [7])) # (!pc_out_2 & ((\btbframes.frameblocks[0].jump_add [7])))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[1].jump_add [7]),
	.datac(\btbframes.frameblocks[0].jump_add [7]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[7]~27_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[7]~27 .lut_mask = 16'hEE50;
defparam \pc_next[7]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N13
dffeas \btbframes.frameblocks[3].jump_add[7] (
	.clk(CLK),
	.d(\pc_when_branch[7]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [7]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[7] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N8
cycloneive_lcell_comb \pc_next[7]~28 (
// Equation(s):
// \pc_next[7]~28_combout  = (pc_out_3 & ((\pc_next[7]~27_combout  & (\btbframes.frameblocks[3].jump_add [7])) # (!\pc_next[7]~27_combout  & ((\btbframes.frameblocks[2].jump_add [7]))))) # (!pc_out_3 & (((\pc_next[7]~27_combout ))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[3].jump_add [7]),
	.datac(\btbframes.frameblocks[2].jump_add [7]),
	.datad(\pc_next[7]~27_combout ),
	.cin(gnd),
	.combout(\pc_next[7]~28_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[7]~28 .lut_mask = 16'hDDA0;
defparam \pc_next[7]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N28
cycloneive_lcell_comb \pc_next[6]~29 (
// Equation(s):
// \pc_next[6]~29_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & ((\pc_when_branch[6]~8_combout ))) # (!pc_out_101 & (pc_plus_4_M[6])))) # (!\branch_or_jump~2_combout  & (pc_out_101))

	.dataa(\branch_or_jump~2_combout ),
	.datab(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datac(pc_plus_4_M[6]),
	.datad(\pc_when_branch[6]~8_combout ),
	.cin(gnd),
	.combout(\pc_next[6]~29_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[6]~29 .lut_mask = 16'hEC64;
defparam \pc_next[6]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N6
cycloneive_lcell_comb \pc_next[6]~30 (
// Equation(s):
// \pc_next[6]~30_combout  = (\branch_or_jump~2_combout  & (((\pc_next[6]~29_combout )))) # (!\branch_or_jump~2_combout  & ((\pc_next[6]~29_combout  & ((imm_M[4]))) # (!\pc_next[6]~29_combout  & (rdata1_M[6]))))

	.dataa(rdata1_M[6]),
	.datab(imm_M[4]),
	.datac(\branch_or_jump~2_combout ),
	.datad(\pc_next[6]~29_combout ),
	.cin(gnd),
	.combout(\pc_next[6]~30_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[6]~30 .lut_mask = 16'hFC0A;
defparam \pc_next[6]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N5
dffeas \btbframes.frameblocks[1].jump_add[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[6]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [6]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[6] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N25
dffeas \btbframes.frameblocks[2].jump_add[6] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [6]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[6] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N19
dffeas \btbframes.frameblocks[0].jump_add[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[6]~8_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [6]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[6] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N18
cycloneive_lcell_comb \pc_next[6]~31 (
// Equation(s):
// \pc_next[6]~31_combout  = (pc_out_2 & (pc_out_3)) # (!pc_out_2 & ((pc_out_3 & ((\btbframes.frameblocks[2].jump_add [6]))) # (!pc_out_3 & (\btbframes.frameblocks[0].jump_add [6]))))

	.dataa(pc_out_2),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[0].jump_add [6]),
	.datad(\btbframes.frameblocks[2].jump_add [6]),
	.cin(gnd),
	.combout(\pc_next[6]~31_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[6]~31 .lut_mask = 16'hDC98;
defparam \pc_next[6]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N11
dffeas \btbframes.frameblocks[3].jump_add[6] (
	.clk(CLK),
	.d(\pc_when_branch[6]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [6]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[6] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N4
cycloneive_lcell_comb \pc_next[6]~32 (
// Equation(s):
// \pc_next[6]~32_combout  = (\pc_next[6]~31_combout  & ((\btbframes.frameblocks[3].jump_add [6]) # ((!pc_out_2)))) # (!\pc_next[6]~31_combout  & (((\btbframes.frameblocks[1].jump_add [6] & pc_out_2))))

	.dataa(\btbframes.frameblocks[3].jump_add [6]),
	.datab(\pc_next[6]~31_combout ),
	.datac(\btbframes.frameblocks[1].jump_add [6]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[6]~32_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[6]~32 .lut_mask = 16'hB8CC;
defparam \pc_next[6]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N24
cycloneive_lcell_comb \pc_next[9]~33 (
// Equation(s):
// \pc_next[9]~33_combout  = (\branch_or_jump~2_combout  & (((pc_plus_4_M[9] & !pc_out_101)))) # (!\branch_or_jump~2_combout  & ((rdata1_M[9]) # ((pc_out_101))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(rdata1_M[9]),
	.datac(pc_plus_4_M[9]),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[9]~33_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[9]~33 .lut_mask = 16'h55E4;
defparam \pc_next[9]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N18
cycloneive_lcell_comb \pc_next[9]~34 (
// Equation(s):
// \pc_next[9]~34_combout  = (pc_out_101 & ((\pc_next[9]~33_combout  & ((imm_M[7]))) # (!\pc_next[9]~33_combout  & (\pc_when_branch[9]~14_combout )))) # (!pc_out_101 & (((\pc_next[9]~33_combout ))))

	.dataa(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datab(\pc_when_branch[9]~14_combout ),
	.datac(imm_M[7]),
	.datad(\pc_next[9]~33_combout ),
	.cin(gnd),
	.combout(\pc_next[9]~34_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[9]~34 .lut_mask = 16'hF588;
defparam \pc_next[9]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N17
dffeas \btbframes.frameblocks[2].jump_add[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[9]~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [9]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[9] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N17
dffeas \btbframes.frameblocks[1].jump_add[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[9]~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [9]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[9] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N31
dffeas \btbframes.frameblocks[0].jump_add[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[9]~14_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [9]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[9] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N30
cycloneive_lcell_comb \pc_next[9]~35 (
// Equation(s):
// \pc_next[9]~35_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].jump_add [9])) # (!pc_out_2 & ((\btbframes.frameblocks[0].jump_add [9])))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[1].jump_add [9]),
	.datac(\btbframes.frameblocks[0].jump_add [9]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[9]~35_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[9]~35 .lut_mask = 16'hEE50;
defparam \pc_next[9]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N17
dffeas \btbframes.frameblocks[3].jump_add[9] (
	.clk(CLK),
	.d(\pc_when_branch[9]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [9]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[9] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N16
cycloneive_lcell_comb \pc_next[9]~36 (
// Equation(s):
// \pc_next[9]~36_combout  = (pc_out_3 & ((\pc_next[9]~35_combout  & ((\btbframes.frameblocks[3].jump_add [9]))) # (!\pc_next[9]~35_combout  & (\btbframes.frameblocks[2].jump_add [9])))) # (!pc_out_3 & (\pc_next[9]~35_combout ))

	.dataa(pc_out_3),
	.datab(\pc_next[9]~35_combout ),
	.datac(\btbframes.frameblocks[2].jump_add [9]),
	.datad(\btbframes.frameblocks[3].jump_add [9]),
	.cin(gnd),
	.combout(\pc_next[9]~36_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[9]~36 .lut_mask = 16'hEC64;
defparam \pc_next[9]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N28
cycloneive_lcell_comb \pc_next[8]~37 (
// Equation(s):
// \pc_next[8]~37_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & ((\pc_when_branch[8]~12_combout ))) # (!pc_out_101 & (pc_plus_4_M[8])))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_M[8]),
	.datac(\pc_when_branch[8]~12_combout ),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[8]~37_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[8]~37 .lut_mask = 16'hF588;
defparam \pc_next[8]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N2
cycloneive_lcell_comb \pc_next[8]~38 (
// Equation(s):
// \pc_next[8]~38_combout  = (\pc_next[8]~37_combout  & (((imm_M[6]) # (\branch_or_jump~2_combout )))) # (!\pc_next[8]~37_combout  & (rdata1_M[8] & ((!\branch_or_jump~2_combout ))))

	.dataa(rdata1_M[8]),
	.datab(\pc_next[8]~37_combout ),
	.datac(imm_M[6]),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\pc_next[8]~38_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[8]~38 .lut_mask = 16'hCCE2;
defparam \pc_next[8]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N25
dffeas \btbframes.frameblocks[1].jump_add[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[8]~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [8]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[8] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N27
dffeas \btbframes.frameblocks[2].jump_add[8] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [8]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[8] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N13
dffeas \btbframes.frameblocks[0].jump_add[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[8]~12_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [8]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[8] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N12
cycloneive_lcell_comb \pc_next[8]~39 (
// Equation(s):
// \pc_next[8]~39_combout  = (pc_out_3 & ((\btbframes.frameblocks[2].jump_add [8]) # ((pc_out_2)))) # (!pc_out_3 & (((\btbframes.frameblocks[0].jump_add [8] & !pc_out_2))))

	.dataa(\btbframes.frameblocks[2].jump_add [8]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[0].jump_add [8]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[8]~39_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[8]~39 .lut_mask = 16'hCCB8;
defparam \pc_next[8]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N15
dffeas \btbframes.frameblocks[3].jump_add[8] (
	.clk(CLK),
	.d(\pc_when_branch[8]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [8]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[8] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N24
cycloneive_lcell_comb \pc_next[8]~40 (
// Equation(s):
// \pc_next[8]~40_combout  = (pc_out_2 & ((\pc_next[8]~39_combout  & ((\btbframes.frameblocks[3].jump_add [8]))) # (!\pc_next[8]~39_combout  & (\btbframes.frameblocks[1].jump_add [8])))) # (!pc_out_2 & (\pc_next[8]~39_combout ))

	.dataa(pc_out_2),
	.datab(\pc_next[8]~39_combout ),
	.datac(\btbframes.frameblocks[1].jump_add [8]),
	.datad(\btbframes.frameblocks[3].jump_add [8]),
	.cin(gnd),
	.combout(\pc_next[8]~40_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[8]~40 .lut_mask = 16'hEC64;
defparam \pc_next[8]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N0
cycloneive_lcell_comb \pc_next[11]~41 (
// Equation(s):
// \pc_next[11]~41_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_M[11] & ((!pc_out_101)))) # (!\branch_or_jump~2_combout  & (((rdata1_M[11]) # (pc_out_101))))

	.dataa(pc_plus_4_M[11]),
	.datab(rdata1_M[11]),
	.datac(\branch_or_jump~2_combout ),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[11]~41_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[11]~41 .lut_mask = 16'h0FAC;
defparam \pc_next[11]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N18
cycloneive_lcell_comb \pc_next[11]~42 (
// Equation(s):
// \pc_next[11]~42_combout  = (pc_out_101 & ((\pc_next[11]~41_combout  & ((imm_M[9]))) # (!\pc_next[11]~41_combout  & (\pc_when_branch[11]~18_combout )))) # (!pc_out_101 & (((\pc_next[11]~41_combout ))))

	.dataa(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datab(\pc_when_branch[11]~18_combout ),
	.datac(imm_M[9]),
	.datad(\pc_next[11]~41_combout ),
	.cin(gnd),
	.combout(\pc_next[11]~42_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[11]~42 .lut_mask = 16'hF588;
defparam \pc_next[11]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N1
dffeas \btbframes.frameblocks[2].jump_add[11] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [11]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[11] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N19
dffeas \btbframes.frameblocks[1].jump_add[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[11]~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [11]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[11] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N29
dffeas \btbframes.frameblocks[0].jump_add[11] (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].jump_add[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [11]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[11] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N18
cycloneive_lcell_comb \pc_next[11]~43 (
// Equation(s):
// \pc_next[11]~43_combout  = (pc_out_2 & ((pc_out_3) # ((\btbframes.frameblocks[1].jump_add [11])))) # (!pc_out_2 & (!pc_out_3 & ((\btbframes.frameblocks[0].jump_add [11]))))

	.dataa(pc_out_2),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[1].jump_add [11]),
	.datad(\btbframes.frameblocks[0].jump_add [11]),
	.cin(gnd),
	.combout(\pc_next[11]~43_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[11]~43 .lut_mask = 16'hB9A8;
defparam \pc_next[11]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N31
dffeas \btbframes.frameblocks[3].jump_add[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[11]~18_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [11]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[11] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N30
cycloneive_lcell_comb \pc_next[11]~44 (
// Equation(s):
// \pc_next[11]~44_combout  = (pc_out_3 & ((\pc_next[11]~43_combout  & ((\btbframes.frameblocks[3].jump_add [11]))) # (!\pc_next[11]~43_combout  & (\btbframes.frameblocks[2].jump_add [11])))) # (!pc_out_3 & (((\pc_next[11]~43_combout ))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[2].jump_add [11]),
	.datac(\btbframes.frameblocks[3].jump_add [11]),
	.datad(\pc_next[11]~43_combout ),
	.cin(gnd),
	.combout(\pc_next[11]~44_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[11]~44 .lut_mask = 16'hF588;
defparam \pc_next[11]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N26
cycloneive_lcell_comb \pc_next[10]~45 (
// Equation(s):
// \pc_next[10]~45_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & ((\pc_when_branch[10]~16_combout ))) # (!pc_out_101 & (pc_plus_4_M[10])))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_M[10]),
	.datac(\pc_when_branch[10]~16_combout ),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[10]~45_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[10]~45 .lut_mask = 16'hF588;
defparam \pc_next[10]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N16
cycloneive_lcell_comb \pc_next[10]~46 (
// Equation(s):
// \pc_next[10]~46_combout  = (\pc_next[10]~45_combout  & ((imm_M[8]) # ((\branch_or_jump~2_combout )))) # (!\pc_next[10]~45_combout  & (((rdata1_M[10] & !\branch_or_jump~2_combout ))))

	.dataa(imm_M[8]),
	.datab(rdata1_M[10]),
	.datac(\pc_next[10]~45_combout ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\pc_next[10]~46_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[10]~46 .lut_mask = 16'hF0AC;
defparam \pc_next[10]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N17
dffeas \btbframes.frameblocks[1].jump_add[10] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[10]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [10]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[10] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N31
dffeas \btbframes.frameblocks[2].jump_add[10] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[10]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [10]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[10] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N21
dffeas \btbframes.frameblocks[0].jump_add[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[10]~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [10]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[10] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N20
cycloneive_lcell_comb \pc_next[10]~47 (
// Equation(s):
// \pc_next[10]~47_combout  = (pc_out_3 & ((\btbframes.frameblocks[2].jump_add [10]) # ((pc_out_2)))) # (!pc_out_3 & (((\btbframes.frameblocks[0].jump_add [10] & !pc_out_2))))

	.dataa(\btbframes.frameblocks[2].jump_add [10]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[0].jump_add [10]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[10]~47_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[10]~47 .lut_mask = 16'hCCB8;
defparam \pc_next[10]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N23
dffeas \btbframes.frameblocks[3].jump_add[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[10]~16_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [10]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[10] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N22
cycloneive_lcell_comb \pc_next[10]~48 (
// Equation(s):
// \pc_next[10]~48_combout  = (pc_out_2 & ((\pc_next[10]~47_combout  & ((\btbframes.frameblocks[3].jump_add [10]))) # (!\pc_next[10]~47_combout  & (\btbframes.frameblocks[1].jump_add [10])))) # (!pc_out_2 & (((\pc_next[10]~47_combout ))))

	.dataa(pc_out_2),
	.datab(\btbframes.frameblocks[1].jump_add [10]),
	.datac(\btbframes.frameblocks[3].jump_add [10]),
	.datad(\pc_next[10]~47_combout ),
	.cin(gnd),
	.combout(\pc_next[10]~48_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[10]~48 .lut_mask = 16'hF588;
defparam \pc_next[10]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N0
cycloneive_lcell_comb \pc_next[13]~49 (
// Equation(s):
// \pc_next[13]~49_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_M[13] & ((!pc_out_101)))) # (!\branch_or_jump~2_combout  & (((rdata1_M[13]) # (pc_out_101))))

	.dataa(pc_plus_4_M[13]),
	.datab(\branch_or_jump~2_combout ),
	.datac(rdata1_M[13]),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[13]~49_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[13]~49 .lut_mask = 16'h33B8;
defparam \pc_next[13]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N18
cycloneive_lcell_comb \pc_next[13]~50 (
// Equation(s):
// \pc_next[13]~50_combout  = (pc_out_101 & ((\pc_next[13]~49_combout  & ((imm_M[11]))) # (!\pc_next[13]~49_combout  & (\pc_when_branch[13]~22_combout )))) # (!pc_out_101 & (((\pc_next[13]~49_combout ))))

	.dataa(\pc_when_branch[13]~22_combout ),
	.datab(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datac(imm_M[11]),
	.datad(\pc_next[13]~49_combout ),
	.cin(gnd),
	.combout(\pc_next[13]~50_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[13]~50 .lut_mask = 16'hF388;
defparam \pc_next[13]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N21
dffeas \btbframes.frameblocks[2].jump_add[13] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[13]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [13]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[13] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N13
dffeas \btbframes.frameblocks[1].jump_add[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[13]~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [13]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[13] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N27
dffeas \btbframes.frameblocks[0].jump_add[13] (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].jump_add[13]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [13]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[13] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N12
cycloneive_lcell_comb \pc_next[13]~51 (
// Equation(s):
// \pc_next[13]~51_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & ((\btbframes.frameblocks[1].jump_add [13]))) # (!pc_out_2 & (\btbframes.frameblocks[0].jump_add [13]))))

	.dataa(\btbframes.frameblocks[0].jump_add [13]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[1].jump_add [13]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[13]~51_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[13]~51 .lut_mask = 16'hFC22;
defparam \pc_next[13]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N31
dffeas \btbframes.frameblocks[3].jump_add[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[13]~22_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [13]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[13] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N30
cycloneive_lcell_comb \pc_next[13]~52 (
// Equation(s):
// \pc_next[13]~52_combout  = (\pc_next[13]~51_combout  & (((\btbframes.frameblocks[3].jump_add [13]) # (!pc_out_3)))) # (!\pc_next[13]~51_combout  & (\btbframes.frameblocks[2].jump_add [13] & ((pc_out_3))))

	.dataa(\pc_next[13]~51_combout ),
	.datab(\btbframes.frameblocks[2].jump_add [13]),
	.datac(\btbframes.frameblocks[3].jump_add [13]),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\pc_next[13]~52_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[13]~52 .lut_mask = 16'hE4AA;
defparam \pc_next[13]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N22
cycloneive_lcell_comb \pc_next[12]~53 (
// Equation(s):
// \pc_next[12]~53_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & ((\pc_when_branch[12]~20_combout ))) # (!pc_out_101 & (pc_plus_4_M[12])))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_M[12]),
	.datac(\pc_when_branch[12]~20_combout ),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[12]~53_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[12]~53 .lut_mask = 16'hF588;
defparam \pc_next[12]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N0
cycloneive_lcell_comb \pc_next[12]~54 (
// Equation(s):
// \pc_next[12]~54_combout  = (\pc_next[12]~53_combout  & (((imm_M[10]) # (\branch_or_jump~2_combout )))) # (!\pc_next[12]~53_combout  & (rdata1_M[12] & ((!\branch_or_jump~2_combout ))))

	.dataa(rdata1_M[12]),
	.datab(imm_M[10]),
	.datac(\pc_next[12]~53_combout ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\pc_next[12]~54_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[12]~54 .lut_mask = 16'hF0CA;
defparam \pc_next[12]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N25
dffeas \btbframes.frameblocks[1].jump_add[12] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[12]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [12]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[12] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N23
dffeas \btbframes.frameblocks[2].jump_add[12] (
	.clk(CLK),
	.d(\pc_when_branch[12]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [12]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[12] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N15
dffeas \btbframes.frameblocks[0].jump_add[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[12]~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [12]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[12] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N14
cycloneive_lcell_comb \pc_next[12]~55 (
// Equation(s):
// \pc_next[12]~55_combout  = (pc_out_3 & ((\btbframes.frameblocks[2].jump_add [12]) # ((pc_out_2)))) # (!pc_out_3 & (((\btbframes.frameblocks[0].jump_add [12] & !pc_out_2))))

	.dataa(\btbframes.frameblocks[2].jump_add [12]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[0].jump_add [12]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[12]~55_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[12]~55 .lut_mask = 16'hCCB8;
defparam \pc_next[12]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N19
dffeas \btbframes.frameblocks[3].jump_add[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[12]~20_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [12]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[12] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N18
cycloneive_lcell_comb \pc_next[12]~56 (
// Equation(s):
// \pc_next[12]~56_combout  = (\pc_next[12]~55_combout  & (((\btbframes.frameblocks[3].jump_add [12]) # (!pc_out_2)))) # (!\pc_next[12]~55_combout  & (\btbframes.frameblocks[1].jump_add [12] & ((pc_out_2))))

	.dataa(\pc_next[12]~55_combout ),
	.datab(\btbframes.frameblocks[1].jump_add [12]),
	.datac(\btbframes.frameblocks[3].jump_add [12]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[12]~56_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[12]~56 .lut_mask = 16'hE4AA;
defparam \pc_next[12]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N8
cycloneive_lcell_comb \pc_next[15]~57 (
// Equation(s):
// \pc_next[15]~57_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_M[15] & ((!pc_out_101)))) # (!\branch_or_jump~2_combout  & (((rdata1_M[15]) # (pc_out_101))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_M[15]),
	.datac(rdata1_M[15]),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[15]~57_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[15]~57 .lut_mask = 16'h55D8;
defparam \pc_next[15]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N16
cycloneive_lcell_comb \pc_next[15]~58 (
// Equation(s):
// \pc_next[15]~58_combout  = (pc_out_101 & ((\pc_next[15]~57_combout  & (imm_M[13])) # (!\pc_next[15]~57_combout  & ((\pc_when_branch[15]~26_combout ))))) # (!pc_out_101 & (((\pc_next[15]~57_combout ))))

	.dataa(imm_M[13]),
	.datab(\pc_when_branch[15]~26_combout ),
	.datac(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datad(\pc_next[15]~57_combout ),
	.cin(gnd),
	.combout(\pc_next[15]~58_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[15]~58 .lut_mask = 16'hAFC0;
defparam \pc_next[15]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y37_N29
dffeas \btbframes.frameblocks[2].jump_add[15] (
	.clk(CLK),
	.d(\pc_when_branch[15]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [15]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[15] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N21
dffeas \btbframes.frameblocks[1].jump_add[15] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [15]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[15] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N25
dffeas \btbframes.frameblocks[0].jump_add[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[15]~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [15]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[15] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N24
cycloneive_lcell_comb \pc_next[15]~59 (
// Equation(s):
// \pc_next[15]~59_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].jump_add [15])) # (!pc_out_2 & ((\btbframes.frameblocks[0].jump_add [15])))))

	.dataa(\btbframes.frameblocks[1].jump_add [15]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[0].jump_add [15]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[15]~59_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[15]~59 .lut_mask = 16'hEE30;
defparam \pc_next[15]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N23
dffeas \btbframes.frameblocks[3].jump_add[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[15]~26_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [15]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[15] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N22
cycloneive_lcell_comb \pc_next[15]~60 (
// Equation(s):
// \pc_next[15]~60_combout  = (pc_out_3 & ((\pc_next[15]~59_combout  & (\btbframes.frameblocks[3].jump_add [15])) # (!\pc_next[15]~59_combout  & ((\btbframes.frameblocks[2].jump_add [15]))))) # (!pc_out_3 & (\pc_next[15]~59_combout ))

	.dataa(pc_out_3),
	.datab(\pc_next[15]~59_combout ),
	.datac(\btbframes.frameblocks[3].jump_add [15]),
	.datad(\btbframes.frameblocks[2].jump_add [15]),
	.cin(gnd),
	.combout(\pc_next[15]~60_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[15]~60 .lut_mask = 16'hE6C4;
defparam \pc_next[15]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N2
cycloneive_lcell_comb \pc_next[14]~61 (
// Equation(s):
// \pc_next[14]~61_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & ((\pc_when_branch[14]~24_combout ))) # (!pc_out_101 & (pc_plus_4_M[14])))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(pc_plus_4_M[14]),
	.datab(\pc_when_branch[14]~24_combout ),
	.datac(\branch_or_jump~2_combout ),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[14]~61_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[14]~61 .lut_mask = 16'hCFA0;
defparam \pc_next[14]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N14
cycloneive_lcell_comb \pc_next[14]~62 (
// Equation(s):
// \pc_next[14]~62_combout  = (\branch_or_jump~2_combout  & (((\pc_next[14]~61_combout )))) # (!\branch_or_jump~2_combout  & ((\pc_next[14]~61_combout  & ((imm_M[12]))) # (!\pc_next[14]~61_combout  & (rdata1_M[14]))))

	.dataa(rdata1_M[14]),
	.datab(imm_M[12]),
	.datac(\branch_or_jump~2_combout ),
	.datad(\pc_next[14]~61_combout ),
	.cin(gnd),
	.combout(\pc_next[14]~62_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[14]~62 .lut_mask = 16'hFC0A;
defparam \pc_next[14]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N25
dffeas \btbframes.frameblocks[1].jump_add[14] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [14]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[14] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N7
dffeas \btbframes.frameblocks[2].jump_add[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[14]~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [14]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[14] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N17
dffeas \btbframes.frameblocks[0].jump_add[14] (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].jump_add[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [14]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[14] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N6
cycloneive_lcell_comb \pc_next[14]~63 (
// Equation(s):
// \pc_next[14]~63_combout  = (pc_out_3 & (((\btbframes.frameblocks[2].jump_add [14]) # (pc_out_2)))) # (!pc_out_3 & (\btbframes.frameblocks[0].jump_add [14] & ((!pc_out_2))))

	.dataa(\btbframes.frameblocks[0].jump_add [14]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[2].jump_add [14]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[14]~63_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[14]~63 .lut_mask = 16'hCCE2;
defparam \pc_next[14]~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N23
dffeas \btbframes.frameblocks[3].jump_add[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[14]~24_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [14]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[14] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N22
cycloneive_lcell_comb \pc_next[14]~64 (
// Equation(s):
// \pc_next[14]~64_combout  = (\pc_next[14]~63_combout  & (((\btbframes.frameblocks[3].jump_add [14])) # (!pc_out_2))) # (!\pc_next[14]~63_combout  & (pc_out_2 & ((\btbframes.frameblocks[1].jump_add [14]))))

	.dataa(\pc_next[14]~63_combout ),
	.datab(pc_out_2),
	.datac(\btbframes.frameblocks[3].jump_add [14]),
	.datad(\btbframes.frameblocks[1].jump_add [14]),
	.cin(gnd),
	.combout(\pc_next[14]~64_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[14]~64 .lut_mask = 16'hE6A2;
defparam \pc_next[14]~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N7
dffeas \pc_plus_4_M[16] (
	.clk(CLK),
	.d(\pc_plus_4_M~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[16]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[16] .is_wysiwyg = "true";
defparam \pc_plus_4_M[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N16
cycloneive_lcell_comb \pc_next[17]~65 (
// Equation(s):
// \pc_next[17]~65_combout  = (pc_out_101 & (((!\branch_or_jump~2_combout )))) # (!pc_out_101 & ((\branch_or_jump~2_combout  & ((pc_plus_4_M[17]))) # (!\branch_or_jump~2_combout  & (rdata1_M[17]))))

	.dataa(rdata1_M[17]),
	.datab(pc_plus_4_M[17]),
	.datac(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\pc_next[17]~65_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[17]~65 .lut_mask = 16'h0CFA;
defparam \pc_next[17]~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N2
cycloneive_lcell_comb \pc_next[17]~66 (
// Equation(s):
// \pc_next[17]~66_combout  = (pc_out_101 & ((\pc_next[17]~65_combout  & ((imm_M[15]))) # (!\pc_next[17]~65_combout  & (\pc_when_branch[17]~30_combout )))) # (!pc_out_101 & (((\pc_next[17]~65_combout ))))

	.dataa(\pc_when_branch[17]~30_combout ),
	.datab(imm_M[15]),
	.datac(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datad(\pc_next[17]~65_combout ),
	.cin(gnd),
	.combout(\pc_next[17]~66_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[17]~66 .lut_mask = 16'hCFA0;
defparam \pc_next[17]~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N23
dffeas \btbframes.frameblocks[2].jump_add[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[17]~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [17]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[17] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N5
dffeas \btbframes.frameblocks[1].jump_add[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[17]~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [17]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[17] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N1
dffeas \btbframes.frameblocks[0].jump_add[17] (
	.clk(CLK),
	.d(\pc_when_branch[17]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [17]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[17] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N4
cycloneive_lcell_comb \pc_next[17]~67 (
// Equation(s):
// \pc_next[17]~67_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & ((\btbframes.frameblocks[1].jump_add [17]))) # (!pc_out_2 & (\btbframes.frameblocks[0].jump_add [17]))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[0].jump_add [17]),
	.datac(\btbframes.frameblocks[1].jump_add [17]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[17]~67_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[17]~67 .lut_mask = 16'hFA44;
defparam \pc_next[17]~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N5
dffeas \btbframes.frameblocks[3].jump_add[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[17]~30_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [17]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[17] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N4
cycloneive_lcell_comb \pc_next[17]~68 (
// Equation(s):
// \pc_next[17]~68_combout  = (pc_out_3 & ((\pc_next[17]~67_combout  & ((\btbframes.frameblocks[3].jump_add [17]))) # (!\pc_next[17]~67_combout  & (\btbframes.frameblocks[2].jump_add [17])))) # (!pc_out_3 & (((\pc_next[17]~67_combout ))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[2].jump_add [17]),
	.datac(\btbframes.frameblocks[3].jump_add [17]),
	.datad(\pc_next[17]~67_combout ),
	.cin(gnd),
	.combout(\pc_next[17]~68_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[17]~68 .lut_mask = 16'hF588;
defparam \pc_next[17]~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N12
cycloneive_lcell_comb \pc_next[16]~69 (
// Equation(s):
// \pc_next[16]~69_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & (\pc_when_branch[16]~28_combout )) # (!pc_out_101 & ((pc_plus_4_M[16]))))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(\pc_when_branch[16]~28_combout ),
	.datab(pc_plus_4_M[16]),
	.datac(\branch_or_jump~2_combout ),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[16]~69_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[16]~69 .lut_mask = 16'hAFC0;
defparam \pc_next[16]~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N10
cycloneive_lcell_comb \pc_next[16]~70 (
// Equation(s):
// \pc_next[16]~70_combout  = (\pc_next[16]~69_combout  & ((imm_M[14]) # ((\branch_or_jump~2_combout )))) # (!\pc_next[16]~69_combout  & (((rdata1_M[16] & !\branch_or_jump~2_combout ))))

	.dataa(\pc_next[16]~69_combout ),
	.datab(imm_M[14]),
	.datac(rdata1_M[16]),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\pc_next[16]~70_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[16]~70 .lut_mask = 16'hAAD8;
defparam \pc_next[16]~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N11
dffeas \btbframes.frameblocks[1].jump_add[16] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [16]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[16] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N9
dffeas \btbframes.frameblocks[2].jump_add[16] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [16]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[16] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N31
dffeas \btbframes.frameblocks[0].jump_add[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[16]~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [16]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[16] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N30
cycloneive_lcell_comb \pc_next[16]~71 (
// Equation(s):
// \pc_next[16]~71_combout  = (pc_out_2 & (((pc_out_3)))) # (!pc_out_2 & ((pc_out_3 & (\btbframes.frameblocks[2].jump_add [16])) # (!pc_out_3 & ((\btbframes.frameblocks[0].jump_add [16])))))

	.dataa(pc_out_2),
	.datab(\btbframes.frameblocks[2].jump_add [16]),
	.datac(\btbframes.frameblocks[0].jump_add [16]),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\pc_next[16]~71_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[16]~71 .lut_mask = 16'hEE50;
defparam \pc_next[16]~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N9
dffeas \btbframes.frameblocks[3].jump_add[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[16]~28_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [16]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[16] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N8
cycloneive_lcell_comb \pc_next[16]~72 (
// Equation(s):
// \pc_next[16]~72_combout  = (\pc_next[16]~71_combout  & (((\btbframes.frameblocks[3].jump_add [16])) # (!pc_out_2))) # (!\pc_next[16]~71_combout  & (pc_out_2 & ((\btbframes.frameblocks[1].jump_add [16]))))

	.dataa(\pc_next[16]~71_combout ),
	.datab(pc_out_2),
	.datac(\btbframes.frameblocks[3].jump_add [16]),
	.datad(\btbframes.frameblocks[1].jump_add [16]),
	.cin(gnd),
	.combout(\pc_next[16]~72_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[16]~72 .lut_mask = 16'hE6A2;
defparam \pc_next[16]~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N1
dffeas \pc_plus_4_M[18] (
	.clk(CLK),
	.d(\pc_plus_4_M~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[18]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[18] .is_wysiwyg = "true";
defparam \pc_plus_4_M[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N18
cycloneive_lcell_comb \pc_next[19]~73 (
// Equation(s):
// \pc_next[19]~73_combout  = (\branch_or_jump~2_combout  & (((!pc_out_101 & pc_plus_4_M[19])))) # (!\branch_or_jump~2_combout  & ((rdata1_M[19]) # ((pc_out_101))))

	.dataa(rdata1_M[19]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datad(pc_plus_4_M[19]),
	.cin(gnd),
	.combout(\pc_next[19]~73_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[19]~73 .lut_mask = 16'h3E32;
defparam \pc_next[19]~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N19
dffeas \instruction_M[17] (
	.clk(CLK),
	.d(\instruction_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_M[17]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_M[17] .is_wysiwyg = "true";
defparam \instruction_M[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N4
cycloneive_lcell_comb \pc_next[19]~74 (
// Equation(s):
// \pc_next[19]~74_combout  = (pc_out_101 & ((\pc_next[19]~73_combout  & ((instruction_M[17]))) # (!\pc_next[19]~73_combout  & (\pc_when_branch[19]~34_combout )))) # (!pc_out_101 & (((\pc_next[19]~73_combout ))))

	.dataa(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datab(\pc_when_branch[19]~34_combout ),
	.datac(instruction_M[17]),
	.datad(\pc_next[19]~73_combout ),
	.cin(gnd),
	.combout(\pc_next[19]~74_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[19]~74 .lut_mask = 16'hF588;
defparam \pc_next[19]~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N19
dffeas \btbframes.frameblocks[2].jump_add[19] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [19]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[19] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N31
dffeas \btbframes.frameblocks[1].jump_add[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[19]~34_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [19]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[19] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N5
dffeas \btbframes.frameblocks[0].jump_add[19] (
	.clk(CLK),
	.d(\pc_when_branch[19]~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [19]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[19] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N30
cycloneive_lcell_comb \pc_next[19]~75 (
// Equation(s):
// \pc_next[19]~75_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & ((\btbframes.frameblocks[1].jump_add [19]))) # (!pc_out_2 & (\btbframes.frameblocks[0].jump_add [19]))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[0].jump_add [19]),
	.datac(\btbframes.frameblocks[1].jump_add [19]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[19]~75_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[19]~75 .lut_mask = 16'hFA44;
defparam \pc_next[19]~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y38_N9
dffeas \btbframes.frameblocks[3].jump_add[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[19]~34_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [19]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[19] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N8
cycloneive_lcell_comb \pc_next[19]~76 (
// Equation(s):
// \pc_next[19]~76_combout  = (\pc_next[19]~75_combout  & (((\btbframes.frameblocks[3].jump_add [19]) # (!pc_out_3)))) # (!\pc_next[19]~75_combout  & (\btbframes.frameblocks[2].jump_add [19] & ((pc_out_3))))

	.dataa(\pc_next[19]~75_combout ),
	.datab(\btbframes.frameblocks[2].jump_add [19]),
	.datac(\btbframes.frameblocks[3].jump_add [19]),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\pc_next[19]~76_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[19]~76 .lut_mask = 16'hE4AA;
defparam \pc_next[19]~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N4
cycloneive_lcell_comb \pc_next[18]~77 (
// Equation(s):
// \pc_next[18]~77_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & ((\pc_when_branch[18]~32_combout ))) # (!pc_out_101 & (pc_plus_4_M[18])))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(pc_plus_4_M[18]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datad(\pc_when_branch[18]~32_combout ),
	.cin(gnd),
	.combout(\pc_next[18]~77_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[18]~77 .lut_mask = 16'hF838;
defparam \pc_next[18]~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y39_N31
dffeas \instruction_M[16] (
	.clk(CLK),
	.d(\instruction_M~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_M[16]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_M[16] .is_wysiwyg = "true";
defparam \instruction_M[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N26
cycloneive_lcell_comb \pc_next[18]~78 (
// Equation(s):
// \pc_next[18]~78_combout  = (\branch_or_jump~2_combout  & (((\pc_next[18]~77_combout )))) # (!\branch_or_jump~2_combout  & ((\pc_next[18]~77_combout  & (instruction_M[16])) # (!\pc_next[18]~77_combout  & ((rdata1_M[18])))))

	.dataa(instruction_M[16]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\pc_next[18]~77_combout ),
	.datad(rdata1_M[18]),
	.cin(gnd),
	.combout(\pc_next[18]~78_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[18]~78 .lut_mask = 16'hE3E0;
defparam \pc_next[18]~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N3
dffeas \btbframes.frameblocks[1].jump_add[18] (
	.clk(CLK),
	.d(\pc_when_branch[18]~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [18]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[18] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N15
dffeas \btbframes.frameblocks[2].jump_add[18] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [18]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[18] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N13
dffeas \btbframes.frameblocks[0].jump_add[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[18]~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [18]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[18] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N12
cycloneive_lcell_comb \pc_next[18]~79 (
// Equation(s):
// \pc_next[18]~79_combout  = (pc_out_3 & ((\btbframes.frameblocks[2].jump_add [18]) # ((pc_out_2)))) # (!pc_out_3 & (((\btbframes.frameblocks[0].jump_add [18] & !pc_out_2))))

	.dataa(\btbframes.frameblocks[2].jump_add [18]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[0].jump_add [18]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[18]~79_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[18]~79 .lut_mask = 16'hCCB8;
defparam \pc_next[18]~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N15
dffeas \btbframes.frameblocks[3].jump_add[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[18]~32_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [18]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[18] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N14
cycloneive_lcell_comb \pc_next[18]~80 (
// Equation(s):
// \pc_next[18]~80_combout  = (\pc_next[18]~79_combout  & (((\btbframes.frameblocks[3].jump_add [18]) # (!pc_out_2)))) # (!\pc_next[18]~79_combout  & (\btbframes.frameblocks[1].jump_add [18] & ((pc_out_2))))

	.dataa(\pc_next[18]~79_combout ),
	.datab(\btbframes.frameblocks[1].jump_add [18]),
	.datac(\btbframes.frameblocks[3].jump_add [18]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[18]~80_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[18]~80 .lut_mask = 16'hE4AA;
defparam \pc_next[18]~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y37_N29
dffeas \pc_plus_4_M[21] (
	.clk(CLK),
	.d(\pc_plus_4_M~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[21]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[21] .is_wysiwyg = "true";
defparam \pc_plus_4_M[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N4
cycloneive_lcell_comb \pc_next[21]~81 (
// Equation(s):
// \pc_next[21]~81_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_M[21] & ((!pc_out_101)))) # (!\branch_or_jump~2_combout  & (((rdata1_M[21]) # (pc_out_101))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_M[21]),
	.datac(rdata1_M[21]),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[21]~81_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[21]~81 .lut_mask = 16'h55D8;
defparam \pc_next[21]~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N27
dffeas \instruction_M[19] (
	.clk(CLK),
	.d(\instruction_M~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_M[19]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_M[19] .is_wysiwyg = "true";
defparam \instruction_M[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N2
cycloneive_lcell_comb \pc_next[21]~82 (
// Equation(s):
// \pc_next[21]~82_combout  = (pc_out_101 & ((\pc_next[21]~81_combout  & (instruction_M[19])) # (!\pc_next[21]~81_combout  & ((\pc_when_branch[21]~38_combout ))))) # (!pc_out_101 & (((\pc_next[21]~81_combout ))))

	.dataa(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datab(instruction_M[19]),
	.datac(\pc_next[21]~81_combout ),
	.datad(\pc_when_branch[21]~38_combout ),
	.cin(gnd),
	.combout(\pc_next[21]~82_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[21]~82 .lut_mask = 16'hDAD0;
defparam \pc_next[21]~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N17
dffeas \btbframes.frameblocks[2].jump_add[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[21]~38_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [21]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[21] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N5
dffeas \btbframes.frameblocks[1].jump_add[21] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [21]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[21] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N11
dffeas \btbframes.frameblocks[0].jump_add[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[21]~38_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [21]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[21] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N10
cycloneive_lcell_comb \pc_next[21]~83 (
// Equation(s):
// \pc_next[21]~83_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].jump_add [21])) # (!pc_out_2 & ((\btbframes.frameblocks[0].jump_add [21])))))

	.dataa(\btbframes.frameblocks[1].jump_add [21]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[0].jump_add [21]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[21]~83_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[21]~83 .lut_mask = 16'hEE30;
defparam \pc_next[21]~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N15
dffeas \btbframes.frameblocks[3].jump_add[21] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].jump_add[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [21]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[21] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N16
cycloneive_lcell_comb \pc_next[21]~84 (
// Equation(s):
// \pc_next[21]~84_combout  = (\pc_next[21]~83_combout  & ((\btbframes.frameblocks[3].jump_add [21]) # ((!pc_out_3)))) # (!\pc_next[21]~83_combout  & (((\btbframes.frameblocks[2].jump_add [21] & pc_out_3))))

	.dataa(\pc_next[21]~83_combout ),
	.datab(\btbframes.frameblocks[3].jump_add [21]),
	.datac(\btbframes.frameblocks[2].jump_add [21]),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\pc_next[21]~84_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[21]~84 .lut_mask = 16'hD8AA;
defparam \pc_next[21]~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N0
cycloneive_lcell_comb \pc_next[20]~85 (
// Equation(s):
// \pc_next[20]~85_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & ((\pc_when_branch[20]~36_combout ))) # (!pc_out_101 & (pc_plus_4_M[20])))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(pc_plus_4_M[20]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datad(\pc_when_branch[20]~36_combout ),
	.cin(gnd),
	.combout(\pc_next[20]~85_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[20]~85 .lut_mask = 16'hF838;
defparam \pc_next[20]~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N31
dffeas \instruction_M[18] (
	.clk(CLK),
	.d(\instruction_M~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_M[18]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_M[18] .is_wysiwyg = "true";
defparam \instruction_M[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N20
cycloneive_lcell_comb \pc_next[20]~86 (
// Equation(s):
// \pc_next[20]~86_combout  = (\branch_or_jump~2_combout  & (((\pc_next[20]~85_combout )))) # (!\branch_or_jump~2_combout  & ((\pc_next[20]~85_combout  & (instruction_M[18])) # (!\pc_next[20]~85_combout  & ((rdata1_M[20])))))

	.dataa(instruction_M[18]),
	.datab(\branch_or_jump~2_combout ),
	.datac(rdata1_M[20]),
	.datad(\pc_next[20]~85_combout ),
	.cin(gnd),
	.combout(\pc_next[20]~86_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[20]~86 .lut_mask = 16'hEE30;
defparam \pc_next[20]~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N7
dffeas \btbframes.frameblocks[1].jump_add[20] (
	.clk(CLK),
	.d(\pc_when_branch[20]~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [20]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[20] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N3
dffeas \btbframes.frameblocks[2].jump_add[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[20]~36_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [20]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[20] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N3
dffeas \btbframes.frameblocks[0].jump_add[20] (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].jump_add[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [20]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[20] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N2
cycloneive_lcell_comb \pc_next[20]~87 (
// Equation(s):
// \pc_next[20]~87_combout  = (pc_out_3 & (((\btbframes.frameblocks[2].jump_add [20]) # (pc_out_2)))) # (!pc_out_3 & (\btbframes.frameblocks[0].jump_add [20] & ((!pc_out_2))))

	.dataa(\btbframes.frameblocks[0].jump_add [20]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[2].jump_add [20]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[20]~87_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[20]~87 .lut_mask = 16'hCCE2;
defparam \pc_next[20]~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N25
dffeas \btbframes.frameblocks[3].jump_add[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[20]~36_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [20]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[20] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N24
cycloneive_lcell_comb \pc_next[20]~88 (
// Equation(s):
// \pc_next[20]~88_combout  = (\pc_next[20]~87_combout  & (((\btbframes.frameblocks[3].jump_add [20])) # (!pc_out_2))) # (!\pc_next[20]~87_combout  & (pc_out_2 & ((\btbframes.frameblocks[1].jump_add [20]))))

	.dataa(\pc_next[20]~87_combout ),
	.datab(pc_out_2),
	.datac(\btbframes.frameblocks[3].jump_add [20]),
	.datad(\btbframes.frameblocks[1].jump_add [20]),
	.cin(gnd),
	.combout(\pc_next[20]~88_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[20]~88 .lut_mask = 16'hE6A2;
defparam \pc_next[20]~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N8
cycloneive_lcell_comb \pc_next[23]~89 (
// Equation(s):
// \pc_next[23]~89_combout  = (pc_out_101 & (((!\branch_or_jump~2_combout )))) # (!pc_out_101 & ((\branch_or_jump~2_combout  & (pc_plus_4_M[23])) # (!\branch_or_jump~2_combout  & ((rdata1_M[23])))))

	.dataa(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datab(pc_plus_4_M[23]),
	.datac(\branch_or_jump~2_combout ),
	.datad(rdata1_M[23]),
	.cin(gnd),
	.combout(\pc_next[23]~89_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[23]~89 .lut_mask = 16'h4F4A;
defparam \pc_next[23]~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N5
dffeas \instruction_M[21] (
	.clk(CLK),
	.d(\instruction_M~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_M[21]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_M[21] .is_wysiwyg = "true";
defparam \instruction_M[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N18
cycloneive_lcell_comb \pc_next[23]~90 (
// Equation(s):
// \pc_next[23]~90_combout  = (pc_out_101 & ((\pc_next[23]~89_combout  & ((instruction_M[21]))) # (!\pc_next[23]~89_combout  & (\pc_when_branch[23]~42_combout )))) # (!pc_out_101 & (\pc_next[23]~89_combout ))

	.dataa(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datab(\pc_next[23]~89_combout ),
	.datac(\pc_when_branch[23]~42_combout ),
	.datad(instruction_M[21]),
	.cin(gnd),
	.combout(\pc_next[23]~90_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[23]~90 .lut_mask = 16'hEC64;
defparam \pc_next[23]~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y39_N29
dffeas \btbframes.frameblocks[2].jump_add[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[23]~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [23]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[23] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y39_N21
dffeas \btbframes.frameblocks[1].jump_add[23] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [23]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[23] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N11
dffeas \btbframes.frameblocks[0].jump_add[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[23]~42_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [23]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[23] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N10
cycloneive_lcell_comb \pc_next[23]~91 (
// Equation(s):
// \pc_next[23]~91_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].jump_add [23])) # (!pc_out_2 & ((\btbframes.frameblocks[0].jump_add [23])))))

	.dataa(\btbframes.frameblocks[1].jump_add [23]),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[0].jump_add [23]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[23]~91_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[23]~91 .lut_mask = 16'hEE30;
defparam \pc_next[23]~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N1
dffeas \btbframes.frameblocks[3].jump_add[23] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].jump_add[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [23]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[23] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N28
cycloneive_lcell_comb \pc_next[23]~92 (
// Equation(s):
// \pc_next[23]~92_combout  = (\pc_next[23]~91_combout  & (((\btbframes.frameblocks[3].jump_add [23])) # (!pc_out_3))) # (!\pc_next[23]~91_combout  & (pc_out_3 & (\btbframes.frameblocks[2].jump_add [23])))

	.dataa(\pc_next[23]~91_combout ),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[2].jump_add [23]),
	.datad(\btbframes.frameblocks[3].jump_add [23]),
	.cin(gnd),
	.combout(\pc_next[23]~92_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[23]~92 .lut_mask = 16'hEA62;
defparam \pc_next[23]~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N16
cycloneive_lcell_comb \pc_next[22]~93 (
// Equation(s):
// \pc_next[22]~93_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & (\pc_when_branch[22]~40_combout )) # (!pc_out_101 & ((pc_plus_4_M[22]))))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(\pc_when_branch[22]~40_combout ),
	.datac(pc_plus_4_M[22]),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[22]~93_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[22]~93 .lut_mask = 16'hDDA0;
defparam \pc_next[22]~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N23
dffeas \instruction_M[20] (
	.clk(CLK),
	.d(\instruction_M~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_M[20]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_M[20] .is_wysiwyg = "true";
defparam \instruction_M[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N24
cycloneive_lcell_comb \pc_next[22]~94 (
// Equation(s):
// \pc_next[22]~94_combout  = (\branch_or_jump~2_combout  & (((\pc_next[22]~93_combout )))) # (!\branch_or_jump~2_combout  & ((\pc_next[22]~93_combout  & ((instruction_M[20]))) # (!\pc_next[22]~93_combout  & (rdata1_M[22]))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(rdata1_M[22]),
	.datac(instruction_M[20]),
	.datad(\pc_next[22]~93_combout ),
	.cin(gnd),
	.combout(\pc_next[22]~94_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[22]~94 .lut_mask = 16'hFA44;
defparam \pc_next[22]~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N31
dffeas \btbframes.frameblocks[1].jump_add[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[22]~40_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [22]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[22] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N15
dffeas \btbframes.frameblocks[2].jump_add[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[22]~40_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [22]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[22] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N11
dffeas \btbframes.frameblocks[0].jump_add[22] (
	.clk(CLK),
	.d(\pc_when_branch[22]~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [22]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[22] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N14
cycloneive_lcell_comb \pc_next[22]~95 (
// Equation(s):
// \pc_next[22]~95_combout  = (pc_out_3 & (((\btbframes.frameblocks[2].jump_add [22]) # (pc_out_2)))) # (!pc_out_3 & (\btbframes.frameblocks[0].jump_add [22] & ((!pc_out_2))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[0].jump_add [22]),
	.datac(\btbframes.frameblocks[2].jump_add [22]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[22]~95_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[22]~95 .lut_mask = 16'hAAE4;
defparam \pc_next[22]~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N11
dffeas \btbframes.frameblocks[3].jump_add[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[22]~40_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [22]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[22] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N10
cycloneive_lcell_comb \pc_next[22]~96 (
// Equation(s):
// \pc_next[22]~96_combout  = (\pc_next[22]~95_combout  & (((\btbframes.frameblocks[3].jump_add [22])) # (!pc_out_2))) # (!\pc_next[22]~95_combout  & (pc_out_2 & ((\btbframes.frameblocks[1].jump_add [22]))))

	.dataa(\pc_next[22]~95_combout ),
	.datab(pc_out_2),
	.datac(\btbframes.frameblocks[3].jump_add [22]),
	.datad(\btbframes.frameblocks[1].jump_add [22]),
	.cin(gnd),
	.combout(\pc_next[22]~96_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[22]~96 .lut_mask = 16'hE6A2;
defparam \pc_next[22]~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N18
cycloneive_lcell_comb \pc_next[25]~97 (
// Equation(s):
// \pc_next[25]~97_combout  = (pc_out_101 & (((!\branch_or_jump~2_combout )))) # (!pc_out_101 & ((\branch_or_jump~2_combout  & (pc_plus_4_M[25])) # (!\branch_or_jump~2_combout  & ((rdata1_M[25])))))

	.dataa(pc_plus_4_M[25]),
	.datab(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datac(\branch_or_jump~2_combout ),
	.datad(rdata1_M[25]),
	.cin(gnd),
	.combout(\pc_next[25]~97_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[25]~97 .lut_mask = 16'h2F2C;
defparam \pc_next[25]~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N13
dffeas \instruction_M[23] (
	.clk(CLK),
	.d(\instruction_M~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_M[23]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_M[23] .is_wysiwyg = "true";
defparam \instruction_M[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N2
cycloneive_lcell_comb \pc_next[25]~98 (
// Equation(s):
// \pc_next[25]~98_combout  = (pc_out_101 & ((\pc_next[25]~97_combout  & (instruction_M[23])) # (!\pc_next[25]~97_combout  & ((\pc_when_branch[25]~46_combout ))))) # (!pc_out_101 & (((\pc_next[25]~97_combout ))))

	.dataa(instruction_M[23]),
	.datab(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datac(\pc_when_branch[25]~46_combout ),
	.datad(\pc_next[25]~97_combout ),
	.cin(gnd),
	.combout(\pc_next[25]~98_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[25]~98 .lut_mask = 16'hBBC0;
defparam \pc_next[25]~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N23
dffeas \btbframes.frameblocks[2].jump_add[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[25]~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [25]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[25] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N19
dffeas \btbframes.frameblocks[1].jump_add[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[25]~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [25]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[25] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N5
dffeas \btbframes.frameblocks[0].jump_add[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[25]~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [25]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[25] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N4
cycloneive_lcell_comb \pc_next[25]~99 (
// Equation(s):
// \pc_next[25]~99_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].jump_add [25])) # (!pc_out_2 & ((\btbframes.frameblocks[0].jump_add [25])))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[1].jump_add [25]),
	.datac(\btbframes.frameblocks[0].jump_add [25]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[25]~99_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[25]~99 .lut_mask = 16'hEE50;
defparam \pc_next[25]~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N17
dffeas \btbframes.frameblocks[3].jump_add[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[25]~46_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [25]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[25] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N16
cycloneive_lcell_comb \pc_next[25]~100 (
// Equation(s):
// \pc_next[25]~100_combout  = (\pc_next[25]~99_combout  & (((\btbframes.frameblocks[3].jump_add [25]) # (!pc_out_3)))) # (!\pc_next[25]~99_combout  & (\btbframes.frameblocks[2].jump_add [25] & ((pc_out_3))))

	.dataa(\pc_next[25]~99_combout ),
	.datab(\btbframes.frameblocks[2].jump_add [25]),
	.datac(\btbframes.frameblocks[3].jump_add [25]),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\pc_next[25]~100_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[25]~100 .lut_mask = 16'hE4AA;
defparam \pc_next[25]~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N16
cycloneive_lcell_comb \pc_next[24]~101 (
// Equation(s):
// \pc_next[24]~101_combout  = (pc_out_101 & (((\pc_when_branch[24]~44_combout ) # (!\branch_or_jump~2_combout )))) # (!pc_out_101 & (pc_plus_4_M[24] & (\branch_or_jump~2_combout )))

	.dataa(pc_plus_4_M[24]),
	.datab(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datac(\branch_or_jump~2_combout ),
	.datad(\pc_when_branch[24]~44_combout ),
	.cin(gnd),
	.combout(\pc_next[24]~101_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[24]~101 .lut_mask = 16'hEC2C;
defparam \pc_next[24]~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N29
dffeas \instruction_M[22] (
	.clk(CLK),
	.d(\instruction_M~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_M[22]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_M[22] .is_wysiwyg = "true";
defparam \instruction_M[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N8
cycloneive_lcell_comb \pc_next[24]~102 (
// Equation(s):
// \pc_next[24]~102_combout  = (\branch_or_jump~2_combout  & (((\pc_next[24]~101_combout )))) # (!\branch_or_jump~2_combout  & ((\pc_next[24]~101_combout  & (instruction_M[22])) # (!\pc_next[24]~101_combout  & ((rdata1_M[24])))))

	.dataa(instruction_M[22]),
	.datab(\branch_or_jump~2_combout ),
	.datac(rdata1_M[24]),
	.datad(\pc_next[24]~101_combout ),
	.cin(gnd),
	.combout(\pc_next[24]~102_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[24]~102 .lut_mask = 16'hEE30;
defparam \pc_next[24]~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N15
dffeas \btbframes.frameblocks[1].jump_add[24] (
	.clk(CLK),
	.d(\pc_when_branch[24]~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [24]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[24] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N17
dffeas \btbframes.frameblocks[2].jump_add[24] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [24]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[24] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y39_N27
dffeas \btbframes.frameblocks[0].jump_add[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[24]~44_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [24]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[24] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N26
cycloneive_lcell_comb \pc_next[24]~103 (
// Equation(s):
// \pc_next[24]~103_combout  = (pc_out_2 & (((pc_out_3)))) # (!pc_out_2 & ((pc_out_3 & (\btbframes.frameblocks[2].jump_add [24])) # (!pc_out_3 & ((\btbframes.frameblocks[0].jump_add [24])))))

	.dataa(pc_out_2),
	.datab(\btbframes.frameblocks[2].jump_add [24]),
	.datac(\btbframes.frameblocks[0].jump_add [24]),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\pc_next[24]~103_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[24]~103 .lut_mask = 16'hEE50;
defparam \pc_next[24]~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N7
dffeas \btbframes.frameblocks[3].jump_add[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[24]~44_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [24]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[24] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N6
cycloneive_lcell_comb \pc_next[24]~104 (
// Equation(s):
// \pc_next[24]~104_combout  = (\pc_next[24]~103_combout  & (((\btbframes.frameblocks[3].jump_add [24]) # (!pc_out_2)))) # (!\pc_next[24]~103_combout  & (\btbframes.frameblocks[1].jump_add [24] & ((pc_out_2))))

	.dataa(\btbframes.frameblocks[1].jump_add [24]),
	.datab(\pc_next[24]~103_combout ),
	.datac(\btbframes.frameblocks[3].jump_add [24]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[24]~104_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[24]~104 .lut_mask = 16'hE2CC;
defparam \pc_next[24]~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N4
cycloneive_lcell_comb \pc_next[27]~105 (
// Equation(s):
// \pc_next[27]~105_combout  = (pc_out_101 & (!\branch_or_jump~2_combout )) # (!pc_out_101 & ((\branch_or_jump~2_combout  & (pc_plus_4_M[27])) # (!\branch_or_jump~2_combout  & ((rdata1_M[27])))))

	.dataa(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datab(\branch_or_jump~2_combout ),
	.datac(pc_plus_4_M[27]),
	.datad(rdata1_M[27]),
	.cin(gnd),
	.combout(\pc_next[27]~105_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[27]~105 .lut_mask = 16'h7362;
defparam \pc_next[27]~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N1
dffeas \instruction_M[25] (
	.clk(CLK),
	.d(\instruction_M~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_M[25]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_M[25] .is_wysiwyg = "true";
defparam \instruction_M[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N22
cycloneive_lcell_comb \pc_next[27]~106 (
// Equation(s):
// \pc_next[27]~106_combout  = (pc_out_101 & ((\pc_next[27]~105_combout  & (instruction_M[25])) # (!\pc_next[27]~105_combout  & ((\pc_when_branch[27]~50_combout ))))) # (!pc_out_101 & (((\pc_next[27]~105_combout ))))

	.dataa(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.datab(instruction_M[25]),
	.datac(\pc_next[27]~105_combout ),
	.datad(\pc_when_branch[27]~50_combout ),
	.cin(gnd),
	.combout(\pc_next[27]~106_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[27]~106 .lut_mask = 16'hDAD0;
defparam \pc_next[27]~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y39_N27
dffeas \btbframes.frameblocks[2].jump_add[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[27]~50_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [27]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[27] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N21
dffeas \btbframes.frameblocks[1].jump_add[27] (
	.clk(CLK),
	.d(\pc_when_branch[27]~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [27]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[27] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y39_N9
dffeas \btbframes.frameblocks[0].jump_add[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[27]~50_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [27]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[27] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N8
cycloneive_lcell_comb \pc_next[27]~107 (
// Equation(s):
// \pc_next[27]~107_combout  = (pc_out_3 & (pc_out_2)) # (!pc_out_3 & ((pc_out_2 & ((\btbframes.frameblocks[1].jump_add [27]))) # (!pc_out_2 & (\btbframes.frameblocks[0].jump_add [27]))))

	.dataa(pc_out_3),
	.datab(pc_out_2),
	.datac(\btbframes.frameblocks[0].jump_add [27]),
	.datad(\btbframes.frameblocks[1].jump_add [27]),
	.cin(gnd),
	.combout(\pc_next[27]~107_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[27]~107 .lut_mask = 16'hDC98;
defparam \pc_next[27]~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y39_N15
dffeas \btbframes.frameblocks[3].jump_add[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[27]~50_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [27]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[27] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N14
cycloneive_lcell_comb \pc_next[27]~108 (
// Equation(s):
// \pc_next[27]~108_combout  = (\pc_next[27]~107_combout  & (((\btbframes.frameblocks[3].jump_add [27]) # (!pc_out_3)))) # (!\pc_next[27]~107_combout  & (\btbframes.frameblocks[2].jump_add [27] & ((pc_out_3))))

	.dataa(\btbframes.frameblocks[2].jump_add [27]),
	.datab(\pc_next[27]~107_combout ),
	.datac(\btbframes.frameblocks[3].jump_add [27]),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\pc_next[27]~108_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[27]~108 .lut_mask = 16'hE2CC;
defparam \pc_next[27]~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N28
cycloneive_lcell_comb \pc_next[26]~109 (
// Equation(s):
// \pc_next[26]~109_combout  = (\branch_or_jump~2_combout  & ((pc_out_101 & ((\pc_when_branch[26]~48_combout ))) # (!pc_out_101 & (pc_plus_4_M[26])))) # (!\branch_or_jump~2_combout  & (((pc_out_101))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_M[26]),
	.datac(\pc_when_branch[26]~48_combout ),
	.datad(\PROGRAM_COUNTER|pc_out[10]~31_combout ),
	.cin(gnd),
	.combout(\pc_next[26]~109_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[26]~109 .lut_mask = 16'hF588;
defparam \pc_next[26]~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N23
dffeas \instruction_M[24] (
	.clk(CLK),
	.d(\instruction_M~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_M[24]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_M[24] .is_wysiwyg = "true";
defparam \instruction_M[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N26
cycloneive_lcell_comb \pc_next[26]~110 (
// Equation(s):
// \pc_next[26]~110_combout  = (\branch_or_jump~2_combout  & (((\pc_next[26]~109_combout )))) # (!\branch_or_jump~2_combout  & ((\pc_next[26]~109_combout  & ((instruction_M[24]))) # (!\pc_next[26]~109_combout  & (rdata1_M[26]))))

	.dataa(rdata1_M[26]),
	.datab(instruction_M[24]),
	.datac(\branch_or_jump~2_combout ),
	.datad(\pc_next[26]~109_combout ),
	.cin(gnd),
	.combout(\pc_next[26]~110_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[26]~110 .lut_mask = 16'hFC0A;
defparam \pc_next[26]~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N15
dffeas \btbframes.frameblocks[1].jump_add[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[26]~48_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [26]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[26] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N1
dffeas \btbframes.frameblocks[2].jump_add[26] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[26]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [26]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[26] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N27
dffeas \btbframes.frameblocks[0].jump_add[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[26]~48_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [26]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[26] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N26
cycloneive_lcell_comb \pc_next[26]~111 (
// Equation(s):
// \pc_next[26]~111_combout  = (pc_out_3 & ((\btbframes.frameblocks[2].jump_add [26]) # ((pc_out_2)))) # (!pc_out_3 & (((\btbframes.frameblocks[0].jump_add [26] & !pc_out_2))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[2].jump_add [26]),
	.datac(\btbframes.frameblocks[0].jump_add [26]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[26]~111_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[26]~111 .lut_mask = 16'hAAD8;
defparam \pc_next[26]~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N29
dffeas \btbframes.frameblocks[3].jump_add[26] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].jump_add[26]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [26]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[26] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N14
cycloneive_lcell_comb \pc_next[26]~112 (
// Equation(s):
// \pc_next[26]~112_combout  = (pc_out_2 & ((\pc_next[26]~111_combout  & (\btbframes.frameblocks[3].jump_add [26])) # (!\pc_next[26]~111_combout  & ((\btbframes.frameblocks[1].jump_add [26]))))) # (!pc_out_2 & (((\pc_next[26]~111_combout ))))

	.dataa(\btbframes.frameblocks[3].jump_add [26]),
	.datab(pc_out_2),
	.datac(\btbframes.frameblocks[1].jump_add [26]),
	.datad(\pc_next[26]~111_combout ),
	.cin(gnd),
	.combout(\pc_next[26]~112_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[26]~112 .lut_mask = 16'hBBC0;
defparam \pc_next[26]~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N29
dffeas \btbframes.frameblocks[2].jump_add[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[29]~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [29]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[29] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N5
dffeas \btbframes.frameblocks[1].jump_add[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[29]~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [29]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[29] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N25
dffeas \btbframes.frameblocks[0].jump_add[29] (
	.clk(CLK),
	.d(\pc_when_branch[29]~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [29]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[29] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N4
cycloneive_lcell_comb \pc_next[29]~113 (
// Equation(s):
// \pc_next[29]~113_combout  = (pc_out_2 & ((pc_out_3) # ((\btbframes.frameblocks[1].jump_add [29])))) # (!pc_out_2 & (!pc_out_3 & ((\btbframes.frameblocks[0].jump_add [29]))))

	.dataa(pc_out_2),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[1].jump_add [29]),
	.datad(\btbframes.frameblocks[0].jump_add [29]),
	.cin(gnd),
	.combout(\pc_next[29]~113_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[29]~113 .lut_mask = 16'hB9A8;
defparam \pc_next[29]~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N3
dffeas \btbframes.frameblocks[3].jump_add[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[29]~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [29]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[29] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N2
cycloneive_lcell_comb \pc_next[29]~114 (
// Equation(s):
// \pc_next[29]~114_combout  = (\pc_next[29]~113_combout  & (((\btbframes.frameblocks[3].jump_add [29]) # (!pc_out_3)))) # (!\pc_next[29]~113_combout  & (\btbframes.frameblocks[2].jump_add [29] & ((pc_out_3))))

	.dataa(\pc_next[29]~113_combout ),
	.datab(\btbframes.frameblocks[2].jump_add [29]),
	.datac(\btbframes.frameblocks[3].jump_add [29]),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\pc_next[29]~114_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[29]~114 .lut_mask = 16'hE4AA;
defparam \pc_next[29]~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N23
dffeas \pc_plus_4_M[28] (
	.clk(CLK),
	.d(\pc_plus_4_M~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[28]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[28] .is_wysiwyg = "true";
defparam \pc_plus_4_M[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N20
cycloneive_lcell_comb \pc_next[29]~115 (
// Equation(s):
// \pc_next[29]~115_combout  = (pc_out_292 & ((\pc_when_branch[29]~54_combout ) # ((pc_out_291)))) # (!pc_out_292 & (((pc_plus_4_M[29] & !pc_out_291))))

	.dataa(\PROGRAM_COUNTER|pc_out[29]~30_combout ),
	.datab(\pc_when_branch[29]~54_combout ),
	.datac(pc_plus_4_M[29]),
	.datad(\PROGRAM_COUNTER|pc_out[29]~29_combout ),
	.cin(gnd),
	.combout(\pc_next[29]~115_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[29]~115 .lut_mask = 16'hAAD8;
defparam \pc_next[29]~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N6
cycloneive_lcell_comb \pc_next[29]~116 (
// Equation(s):
// \pc_next[29]~116_combout  = (pc_out_291 & ((\pc_next[29]~115_combout  & (rdata1_M[29])) # (!\pc_next[29]~115_combout  & ((\pc_plus_4[29]~54_combout ))))) # (!pc_out_291 & (((\pc_next[29]~115_combout ))))

	.dataa(\PROGRAM_COUNTER|pc_out[29]~29_combout ),
	.datab(rdata1_M[29]),
	.datac(\pc_plus_4[29]~54_combout ),
	.datad(\pc_next[29]~115_combout ),
	.cin(gnd),
	.combout(\pc_next[29]~116_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[29]~116 .lut_mask = 16'hDDA0;
defparam \pc_next[29]~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N4
cycloneive_lcell_comb \pc_next[29]~117 (
// Equation(s):
// \pc_next[29]~117_combout  = (predicted & ((\branch_or_jump~1_combout  & (\pc_next[29]~114_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[29]~116_combout ))))) # (!predicted & (((\pc_next[29]~116_combout ))))

	.dataa(\BTB|predicted~18_combout ),
	.datab(\pc_next[29]~114_combout ),
	.datac(\branch_or_jump~1_combout ),
	.datad(\pc_next[29]~116_combout ),
	.cin(gnd),
	.combout(\pc_next[29]~117_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[29]~117 .lut_mask = 16'hDF80;
defparam \pc_next[29]~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N31
dffeas \btbframes.frameblocks[1].jump_add[28] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].jump_add[28]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [28]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[28] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N17
dffeas \btbframes.frameblocks[2].jump_add[28] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[28]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [28]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[28] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N3
dffeas \btbframes.frameblocks[0].jump_add[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[28]~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [28]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[28] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N2
cycloneive_lcell_comb \pc_next[28]~118 (
// Equation(s):
// \pc_next[28]~118_combout  = (pc_out_3 & ((\btbframes.frameblocks[2].jump_add [28]) # ((pc_out_2)))) # (!pc_out_3 & (((\btbframes.frameblocks[0].jump_add [28] & !pc_out_2))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[2].jump_add [28]),
	.datac(\btbframes.frameblocks[0].jump_add [28]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[28]~118_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[28]~118 .lut_mask = 16'hAAD8;
defparam \pc_next[28]~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N17
dffeas \btbframes.frameblocks[3].jump_add[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[28]~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [28]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[28] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N16
cycloneive_lcell_comb \pc_next[28]~119 (
// Equation(s):
// \pc_next[28]~119_combout  = (pc_out_2 & ((\pc_next[28]~118_combout  & (\btbframes.frameblocks[3].jump_add [28])) # (!\pc_next[28]~118_combout  & ((\btbframes.frameblocks[1].jump_add [28]))))) # (!pc_out_2 & (\pc_next[28]~118_combout ))

	.dataa(pc_out_2),
	.datab(\pc_next[28]~118_combout ),
	.datac(\btbframes.frameblocks[3].jump_add [28]),
	.datad(\btbframes.frameblocks[1].jump_add [28]),
	.cin(gnd),
	.combout(\pc_next[28]~119_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[28]~119 .lut_mask = 16'hE6C4;
defparam \pc_next[28]~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N28
cycloneive_lcell_comb \pc_next[28]~120 (
// Equation(s):
// \pc_next[28]~120_combout  = (pc_out_292 & (((pc_out_291)))) # (!pc_out_292 & ((pc_out_291 & (\pc_plus_4[28]~52_combout )) # (!pc_out_291 & ((pc_plus_4_M[28])))))

	.dataa(\PROGRAM_COUNTER|pc_out[29]~30_combout ),
	.datab(\pc_plus_4[28]~52_combout ),
	.datac(pc_plus_4_M[28]),
	.datad(\PROGRAM_COUNTER|pc_out[29]~29_combout ),
	.cin(gnd),
	.combout(\pc_next[28]~120_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[28]~120 .lut_mask = 16'hEE50;
defparam \pc_next[28]~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N26
cycloneive_lcell_comb \pc_next[28]~121 (
// Equation(s):
// \pc_next[28]~121_combout  = (pc_out_292 & ((\pc_next[28]~120_combout  & (rdata1_M[28])) # (!\pc_next[28]~120_combout  & ((\pc_when_branch[28]~52_combout ))))) # (!pc_out_292 & (((\pc_next[28]~120_combout ))))

	.dataa(rdata1_M[28]),
	.datab(\PROGRAM_COUNTER|pc_out[29]~30_combout ),
	.datac(\pc_when_branch[28]~52_combout ),
	.datad(\pc_next[28]~120_combout ),
	.cin(gnd),
	.combout(\pc_next[28]~121_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[28]~121 .lut_mask = 16'hBBC0;
defparam \pc_next[28]~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N22
cycloneive_lcell_comb \pc_next[28]~122 (
// Equation(s):
// \pc_next[28]~122_combout  = (\branch_or_jump~1_combout  & ((predicted & ((\pc_next[28]~119_combout ))) # (!predicted & (\pc_next[28]~121_combout )))) # (!\branch_or_jump~1_combout  & (\pc_next[28]~121_combout ))

	.dataa(\pc_next[28]~121_combout ),
	.datab(\pc_next[28]~119_combout ),
	.datac(\branch_or_jump~1_combout ),
	.datad(\BTB|predicted~18_combout ),
	.cin(gnd),
	.combout(\pc_next[28]~122_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[28]~122 .lut_mask = 16'hCAAA;
defparam \pc_next[28]~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N15
dffeas \btbframes.frameblocks[2].jump_add[31] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[31]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [31]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[31] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N29
dffeas \btbframes.frameblocks[1].jump_add[31] (
	.clk(CLK),
	.d(\pc_when_branch[31]~58_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [31]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[31] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N7
dffeas \btbframes.frameblocks[0].jump_add[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[31]~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [31]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[31] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N6
cycloneive_lcell_comb \pc_next[31]~123 (
// Equation(s):
// \pc_next[31]~123_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].jump_add [31])) # (!pc_out_2 & ((\btbframes.frameblocks[0].jump_add [31])))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[1].jump_add [31]),
	.datac(\btbframes.frameblocks[0].jump_add [31]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[31]~123_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[31]~123 .lut_mask = 16'hEE50;
defparam \pc_next[31]~123 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N9
dffeas \btbframes.frameblocks[3].jump_add[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[31]~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [31]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[31] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N8
cycloneive_lcell_comb \pc_next[31]~124 (
// Equation(s):
// \pc_next[31]~124_combout  = (\pc_next[31]~123_combout  & (((\btbframes.frameblocks[3].jump_add [31])) # (!pc_out_3))) # (!\pc_next[31]~123_combout  & (pc_out_3 & ((\btbframes.frameblocks[2].jump_add [31]))))

	.dataa(\pc_next[31]~123_combout ),
	.datab(pc_out_3),
	.datac(\btbframes.frameblocks[3].jump_add [31]),
	.datad(\btbframes.frameblocks[2].jump_add [31]),
	.cin(gnd),
	.combout(\pc_next[31]~124_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[31]~124 .lut_mask = 16'hE6A2;
defparam \pc_next[31]~124 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N12
cycloneive_lcell_comb \pc_next[31]~125 (
// Equation(s):
// \pc_next[31]~125_combout  = (pc_out_291 & (pc_out_292)) # (!pc_out_291 & ((pc_out_292 & ((\pc_when_branch[31]~58_combout ))) # (!pc_out_292 & (pc_plus_4_M[31]))))

	.dataa(\PROGRAM_COUNTER|pc_out[29]~29_combout ),
	.datab(\PROGRAM_COUNTER|pc_out[29]~30_combout ),
	.datac(pc_plus_4_M[31]),
	.datad(\pc_when_branch[31]~58_combout ),
	.cin(gnd),
	.combout(\pc_next[31]~125_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[31]~125 .lut_mask = 16'hDC98;
defparam \pc_next[31]~125 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N30
cycloneive_lcell_comb \pc_next[31]~126 (
// Equation(s):
// \pc_next[31]~126_combout  = (pc_out_291 & ((\pc_next[31]~125_combout  & (rdata1_M[31])) # (!\pc_next[31]~125_combout  & ((\pc_plus_4[31]~58_combout ))))) # (!pc_out_291 & (((\pc_next[31]~125_combout ))))

	.dataa(\PROGRAM_COUNTER|pc_out[29]~29_combout ),
	.datab(rdata1_M[31]),
	.datac(\pc_plus_4[31]~58_combout ),
	.datad(\pc_next[31]~125_combout ),
	.cin(gnd),
	.combout(\pc_next[31]~126_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[31]~126 .lut_mask = 16'hDDA0;
defparam \pc_next[31]~126 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N0
cycloneive_lcell_comb \pc_next[31]~127 (
// Equation(s):
// \pc_next[31]~127_combout  = (\branch_or_jump~1_combout  & ((predicted & (\pc_next[31]~124_combout )) # (!predicted & ((\pc_next[31]~126_combout ))))) # (!\branch_or_jump~1_combout  & (((\pc_next[31]~126_combout ))))

	.dataa(\pc_next[31]~124_combout ),
	.datab(\branch_or_jump~1_combout ),
	.datac(\pc_next[31]~126_combout ),
	.datad(\BTB|predicted~18_combout ),
	.cin(gnd),
	.combout(\pc_next[31]~127_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[31]~127 .lut_mask = 16'hB8F0;
defparam \pc_next[31]~127 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N27
dffeas \btbframes.frameblocks[1].jump_add[30] (
	.clk(CLK),
	.d(\pc_when_branch[30]~56_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].jump_add [30]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[30] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].jump_add[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N13
dffeas \btbframes.frameblocks[2].jump_add[30] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].jump_add[30]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].jump_add [30]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[30] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].jump_add[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N19
dffeas \btbframes.frameblocks[0].jump_add[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[30]~56_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].jump_add [30]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[30] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].jump_add[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N18
cycloneive_lcell_comb \pc_next[30]~128 (
// Equation(s):
// \pc_next[30]~128_combout  = (pc_out_3 & ((\btbframes.frameblocks[2].jump_add [30]) # ((pc_out_2)))) # (!pc_out_3 & (((\btbframes.frameblocks[0].jump_add [30] & !pc_out_2))))

	.dataa(pc_out_3),
	.datab(\btbframes.frameblocks[2].jump_add [30]),
	.datac(\btbframes.frameblocks[0].jump_add [30]),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\pc_next[30]~128_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[30]~128 .lut_mask = 16'hAAD8;
defparam \pc_next[30]~128 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N21
dffeas \btbframes.frameblocks[3].jump_add[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_when_branch[30]~56_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].jump_add [30]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[30] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].jump_add[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N20
cycloneive_lcell_comb \pc_next[30]~129 (
// Equation(s):
// \pc_next[30]~129_combout  = (pc_out_2 & ((\pc_next[30]~128_combout  & (\btbframes.frameblocks[3].jump_add [30])) # (!\pc_next[30]~128_combout  & ((\btbframes.frameblocks[1].jump_add [30]))))) # (!pc_out_2 & (\pc_next[30]~128_combout ))

	.dataa(pc_out_2),
	.datab(\pc_next[30]~128_combout ),
	.datac(\btbframes.frameblocks[3].jump_add [30]),
	.datad(\btbframes.frameblocks[1].jump_add [30]),
	.cin(gnd),
	.combout(\pc_next[30]~129_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[30]~129 .lut_mask = 16'hE6C4;
defparam \pc_next[30]~129 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N30
cycloneive_lcell_comb \pc_next[30]~130 (
// Equation(s):
// \pc_next[30]~130_combout  = (pc_out_291 & ((\pc_plus_4[30]~56_combout ) # ((pc_out_292)))) # (!pc_out_291 & (((pc_plus_4_M[30] & !pc_out_292))))

	.dataa(\PROGRAM_COUNTER|pc_out[29]~29_combout ),
	.datab(\pc_plus_4[30]~56_combout ),
	.datac(pc_plus_4_M[30]),
	.datad(\PROGRAM_COUNTER|pc_out[29]~30_combout ),
	.cin(gnd),
	.combout(\pc_next[30]~130_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[30]~130 .lut_mask = 16'hAAD8;
defparam \pc_next[30]~130 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N0
cycloneive_lcell_comb \pc_next[30]~131 (
// Equation(s):
// \pc_next[30]~131_combout  = (pc_out_292 & ((\pc_next[30]~130_combout  & ((rdata1_M[30]))) # (!\pc_next[30]~130_combout  & (\pc_when_branch[30]~56_combout )))) # (!pc_out_292 & (((\pc_next[30]~130_combout ))))

	.dataa(\PROGRAM_COUNTER|pc_out[29]~30_combout ),
	.datab(\pc_when_branch[30]~56_combout ),
	.datac(\pc_next[30]~130_combout ),
	.datad(rdata1_M[30]),
	.cin(gnd),
	.combout(\pc_next[30]~131_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[30]~131 .lut_mask = 16'hF858;
defparam \pc_next[30]~131 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N14
cycloneive_lcell_comb \pc_next[30]~132 (
// Equation(s):
// \pc_next[30]~132_combout  = (\branch_or_jump~1_combout  & ((predicted & (\pc_next[30]~129_combout )) # (!predicted & ((\pc_next[30]~131_combout ))))) # (!\branch_or_jump~1_combout  & (((\pc_next[30]~131_combout ))))

	.dataa(\pc_next[30]~129_combout ),
	.datab(\branch_or_jump~1_combout ),
	.datac(\pc_next[30]~131_combout ),
	.datad(\BTB|predicted~18_combout ),
	.cin(gnd),
	.combout(\pc_next[30]~132_combout ),
	.cout());
// synopsys translate_off
defparam \pc_next[30]~132 .lut_mask = 16'hB8F0;
defparam \pc_next[30]~132 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N13
dffeas cu_halt_EX(
	.clk(CLK),
	.d(\cu_halt_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\cu_halt_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam cu_halt_EX.is_wysiwyg = "true";
defparam cu_halt_EX.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N21
dffeas jal_EX(
	.clk(CLK),
	.d(\jal_EX~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\jal_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam jal_EX.is_wysiwyg = "true";
defparam jal_EX.power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N25
dffeas predicted_EX(
	.clk(CLK),
	.d(\predicted_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\predicted_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam predicted_EX.is_wysiwyg = "true";
defparam predicted_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N0
cycloneive_lcell_comb \bne_M~0 (
// Equation(s):
// \bne_M~0_combout  = (\bne_EX~q  & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\bne_EX~q ),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\bne_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \bne_M~0 .lut_mask = 16'h00F0;
defparam \bne_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N10
cycloneive_lcell_comb \zero_M~5 (
// Equation(s):
// \zero_M~5_combout  = (Selector30) # ((Selector161) # ((Selector12 & ShiftRight0)))

	.dataa(\ALU|Selector12~10_combout ),
	.datab(\ALU|ShiftRight0~91_combout ),
	.datac(\ALU|Selector30~8_combout ),
	.datad(\ALU|Selector16~11_combout ),
	.cin(gnd),
	.combout(\zero_M~5_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~5 .lut_mask = 16'hFFF8;
defparam \zero_M~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N17
dffeas jr_EX(
	.clk(CLK),
	.d(\jr_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\jr_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam jr_EX.is_wysiwyg = "true";
defparam jr_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N6
cycloneive_lcell_comb \jr_M~0 (
// Equation(s):
// \jr_M~0_combout  = (\jr_EX~q  & (!\en_EX~0_combout  & !\wsel_M~0_combout ))

	.dataa(gnd),
	.datab(\jr_EX~q ),
	.datac(\en_EX~0_combout ),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\jr_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \jr_M~0 .lut_mask = 16'h000C;
defparam \jr_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N5
dffeas \op_D[5] (
	.clk(CLK),
	.d(\op_D~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_D[5]),
	.prn(vcc));
// synopsys translate_off
defparam \op_D[5] .is_wysiwyg = "true";
defparam \op_D[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N8
cycloneive_lcell_comb \op_EX~0 (
// Equation(s):
// \op_EX~0_combout  = ((op_D[5]) # (\predicted_M~q  $ (\branch_taken~0_combout ))) # (!\branch_or_jump~2_combout )

	.dataa(\branch_or_jump~2_combout ),
	.datab(op_D[5]),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\op_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \op_EX~0 .lut_mask = 16'hDFFD;
defparam \op_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N29
dffeas \op_D[4] (
	.clk(CLK),
	.d(\op_D~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_D[4]),
	.prn(vcc));
// synopsys translate_off
defparam \op_D[4] .is_wysiwyg = "true";
defparam \op_D[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N10
cycloneive_lcell_comb \op_EX~1 (
// Equation(s):
// \op_EX~1_combout  = ((op_D[4]) # (\predicted_M~q  $ (\branch_taken~0_combout ))) # (!\branch_or_jump~2_combout )

	.dataa(\predicted_M~q ),
	.datab(\branch_or_jump~2_combout ),
	.datac(op_D[4]),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\op_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \op_EX~1 .lut_mask = 16'hF7FB;
defparam \op_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N15
dffeas \op_D[3] (
	.clk(CLK),
	.d(\op_D~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_D[3]),
	.prn(vcc));
// synopsys translate_off
defparam \op_D[3] .is_wysiwyg = "true";
defparam \op_D[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N16
cycloneive_lcell_comb \op_EX~2 (
// Equation(s):
// \op_EX~2_combout  = ((op_D[3]) # (\predicted_M~q  $ (\branch_taken~0_combout ))) # (!\branch_or_jump~2_combout )

	.dataa(\predicted_M~q ),
	.datab(\branch_or_jump~2_combout ),
	.datac(op_D[3]),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\op_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \op_EX~2 .lut_mask = 16'hF7FB;
defparam \op_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N27
dffeas \op_D[2] (
	.clk(CLK),
	.d(\op_D~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_D[2]),
	.prn(vcc));
// synopsys translate_off
defparam \op_D[2] .is_wysiwyg = "true";
defparam \op_D[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N24
cycloneive_lcell_comb \op_EX~3 (
// Equation(s):
// \op_EX~3_combout  = (op_D[2]) # ((\branch_taken~0_combout  $ (\predicted_M~q )) # (!\branch_or_jump~2_combout ))

	.dataa(op_D[2]),
	.datab(\branch_taken~0_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\op_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \op_EX~3 .lut_mask = 16'hBEFF;
defparam \op_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N9
dffeas \op_D[1] (
	.clk(CLK),
	.d(\op_D~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_D[1]),
	.prn(vcc));
// synopsys translate_off
defparam \op_D[1] .is_wysiwyg = "true";
defparam \op_D[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N22
cycloneive_lcell_comb \op_EX~4 (
// Equation(s):
// \op_EX~4_combout  = ((op_D[1]) # (\predicted_M~q  $ (\branch_taken~0_combout ))) # (!\branch_or_jump~2_combout )

	.dataa(\branch_or_jump~2_combout ),
	.datab(\predicted_M~q ),
	.datac(op_D[1]),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\op_EX~4_combout ),
	.cout());
// synopsys translate_off
defparam \op_EX~4 .lut_mask = 16'hF7FD;
defparam \op_EX~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N7
dffeas \op_D[0] (
	.clk(CLK),
	.d(\op_D~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(op_D[0]),
	.prn(vcc));
// synopsys translate_off
defparam \op_D[0] .is_wysiwyg = "true";
defparam \op_D[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N0
cycloneive_lcell_comb \op_EX~5 (
// Equation(s):
// \op_EX~5_combout  = ((op_D[0]) # (\branch_taken~0_combout  $ (\predicted_M~q ))) # (!\branch_or_jump~2_combout )

	.dataa(\branch_taken~0_combout ),
	.datab(\predicted_M~q ),
	.datac(\branch_or_jump~2_combout ),
	.datad(op_D[0]),
	.cin(gnd),
	.combout(\op_EX~5_combout ),
	.cout());
// synopsys translate_off
defparam \op_EX~5 .lut_mask = 16'hFF6F;
defparam \op_EX~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N29
dffeas \instruction_D[16] (
	.clk(CLK),
	.d(\instruction_D~70_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[16]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[16] .is_wysiwyg = "true";
defparam \instruction_D[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N16
cycloneive_lcell_comb \instruction_EX~0 (
// Equation(s):
// \instruction_EX~0_combout  = (instruction_D[16] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_taken~0_combout ),
	.datab(instruction_D[16]),
	.datac(\predicted_M~q ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\instruction_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_EX~0 .lut_mask = 16'h8400;
defparam \instruction_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N1
dffeas \instruction_D[17] (
	.clk(CLK),
	.d(\instruction_D~71_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[17]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[17] .is_wysiwyg = "true";
defparam \instruction_D[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N30
cycloneive_lcell_comb \instruction_EX~1 (
// Equation(s):
// \instruction_EX~1_combout  = (instruction_D[17] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_taken~0_combout ),
	.datab(instruction_D[17]),
	.datac(\predicted_M~q ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\instruction_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_EX~1 .lut_mask = 16'h8400;
defparam \instruction_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N27
dffeas RegDst_EX(
	.clk(CLK),
	.d(\RegDst_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\RegDst_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam RegDst_EX.is_wysiwyg = "true";
defparam RegDst_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N10
cycloneive_lcell_comb \wsel_M~1 (
// Equation(s):
// \wsel_M~1_combout  = (\RegDst_EX~q  & ((imm_EX[12]))) # (!\RegDst_EX~q  & (instruction_EX[17]))

	.dataa(instruction_EX[17]),
	.datab(gnd),
	.datac(imm_EX[12]),
	.datad(\RegDst_EX~q ),
	.cin(gnd),
	.combout(\wsel_M~1_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~1 .lut_mask = 16'hF0AA;
defparam \wsel_M~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N8
cycloneive_lcell_comb \wsel_M~2 (
// Equation(s):
// \wsel_M~2_combout  = (!\wsel_M~0_combout  & ((\jal_EX~q ) # (\wsel_M~1_combout )))

	.dataa(\wsel_M~0_combout ),
	.datab(gnd),
	.datac(\jal_EX~q ),
	.datad(\wsel_M~1_combout ),
	.cin(gnd),
	.combout(\wsel_M~2_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~2 .lut_mask = 16'h5550;
defparam \wsel_M~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N24
cycloneive_lcell_comb \wsel_M~3 (
// Equation(s):
// \wsel_M~3_combout  = (\RegDst_EX~q  & (imm_EX[11])) # (!\RegDst_EX~q  & ((instruction_EX[16])))

	.dataa(imm_EX[11]),
	.datab(\RegDst_EX~q ),
	.datac(gnd),
	.datad(instruction_EX[16]),
	.cin(gnd),
	.combout(\wsel_M~3_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~3 .lut_mask = 16'hBB88;
defparam \wsel_M~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N2
cycloneive_lcell_comb \wsel_M~4 (
// Equation(s):
// \wsel_M~4_combout  = (!\wsel_M~0_combout  & ((\jal_EX~q ) # (\wsel_M~3_combout )))

	.dataa(\wsel_M~0_combout ),
	.datab(\jal_EX~q ),
	.datac(gnd),
	.datad(\wsel_M~3_combout ),
	.cin(gnd),
	.combout(\wsel_M~4_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~4 .lut_mask = 16'h5544;
defparam \wsel_M~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N7
dffeas \instruction_D[18] (
	.clk(CLK),
	.d(\instruction_D~72_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[18]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[18] .is_wysiwyg = "true";
defparam \instruction_D[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N14
cycloneive_lcell_comb \instruction_EX~2 (
// Equation(s):
// \instruction_EX~2_combout  = (instruction_D[18] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_taken~0_combout ),
	.datab(instruction_D[18]),
	.datac(\predicted_M~q ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\instruction_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_EX~2 .lut_mask = 16'h8400;
defparam \instruction_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N31
dffeas \instruction_D[19] (
	.clk(CLK),
	.d(\instruction_D~73_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[19]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[19] .is_wysiwyg = "true";
defparam \instruction_D[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N28
cycloneive_lcell_comb \instruction_EX~3 (
// Equation(s):
// \instruction_EX~3_combout  = (\branch_or_jump~2_combout  & (instruction_D[19] & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(instruction_D[19]),
	.datac(\branch_taken~0_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\instruction_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_EX~3 .lut_mask = 16'h8008;
defparam \instruction_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N24
cycloneive_lcell_comb \wsel_M~5 (
// Equation(s):
// \wsel_M~5_combout  = (\RegDst_EX~q  & ((imm_EX[14]))) # (!\RegDst_EX~q  & (instruction_EX[19]))

	.dataa(instruction_EX[19]),
	.datab(imm_EX[14]),
	.datac(gnd),
	.datad(\RegDst_EX~q ),
	.cin(gnd),
	.combout(\wsel_M~5_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~5 .lut_mask = 16'hCCAA;
defparam \wsel_M~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N26
cycloneive_lcell_comb \wsel_M~6 (
// Equation(s):
// \wsel_M~6_combout  = (!\wsel_M~0_combout  & ((\jal_EX~q ) # (\wsel_M~5_combout )))

	.dataa(gnd),
	.datab(\jal_EX~q ),
	.datac(\wsel_M~5_combout ),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\wsel_M~6_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~6 .lut_mask = 16'h00FC;
defparam \wsel_M~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N28
cycloneive_lcell_comb \wsel_M~7 (
// Equation(s):
// \wsel_M~7_combout  = (\RegDst_EX~q  & ((imm_EX[13]))) # (!\RegDst_EX~q  & (instruction_EX[18]))

	.dataa(gnd),
	.datab(instruction_EX[18]),
	.datac(\RegDst_EX~q ),
	.datad(imm_EX[13]),
	.cin(gnd),
	.combout(\wsel_M~7_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~7 .lut_mask = 16'hFC0C;
defparam \wsel_M~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N4
cycloneive_lcell_comb \wsel_M~8 (
// Equation(s):
// \wsel_M~8_combout  = (!\wsel_M~0_combout  & ((\jal_EX~q ) # (\wsel_M~7_combout )))

	.dataa(\wsel_M~0_combout ),
	.datab(\jal_EX~q ),
	.datac(gnd),
	.datad(\wsel_M~7_combout ),
	.cin(gnd),
	.combout(\wsel_M~8_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~8 .lut_mask = 16'h5544;
defparam \wsel_M~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N14
cycloneive_lcell_comb \instruction_EX~4 (
// Equation(s):
// \instruction_EX~4_combout  = (instruction_D[20] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(instruction_D[20]),
	.datab(\branch_taken~0_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\instruction_EX~4_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_EX~4 .lut_mask = 16'h8200;
defparam \instruction_EX~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N16
cycloneive_lcell_comb \wsel_M~9 (
// Equation(s):
// \wsel_M~9_combout  = (\RegDst_EX~q  & (imm_EX[15])) # (!\RegDst_EX~q  & ((instruction_EX[20])))

	.dataa(gnd),
	.datab(imm_EX[15]),
	.datac(instruction_EX[20]),
	.datad(\RegDst_EX~q ),
	.cin(gnd),
	.combout(\wsel_M~9_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~9 .lut_mask = 16'hCCF0;
defparam \wsel_M~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N20
cycloneive_lcell_comb \wsel_M~10 (
// Equation(s):
// \wsel_M~10_combout  = (!\wsel_M~0_combout  & ((\wsel_M~9_combout ) # (\jal_EX~q )))

	.dataa(\wsel_M~0_combout ),
	.datab(\wsel_M~9_combout ),
	.datac(\jal_EX~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\wsel_M~10_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~10 .lut_mask = 16'h5454;
defparam \wsel_M~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N9
dffeas \instruction_D[22] (
	.clk(CLK),
	.d(\instruction_D~75_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[22]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[22] .is_wysiwyg = "true";
defparam \instruction_D[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N6
cycloneive_lcell_comb \instruction_EX~5 (
// Equation(s):
// \instruction_EX~5_combout  = (instruction_D[22] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(instruction_D[22]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\branch_taken~0_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\instruction_EX~5_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_EX~5 .lut_mask = 16'h8008;
defparam \instruction_EX~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N9
dffeas \instruction_D[24] (
	.clk(CLK),
	.d(\instruction_D~77_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[24]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[24] .is_wysiwyg = "true";
defparam \instruction_D[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N0
cycloneive_lcell_comb \instruction_EX~7 (
// Equation(s):
// \instruction_EX~7_combout  = (\branch_or_jump~2_combout  & (instruction_D[24] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(\branch_or_jump~2_combout ),
	.datac(\branch_taken~0_combout ),
	.datad(instruction_D[24]),
	.cin(gnd),
	.combout(\instruction_EX~7_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_EX~7 .lut_mask = 16'h8400;
defparam \instruction_EX~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N15
dffeas \instruction_D[23] (
	.clk(CLK),
	.d(\instruction_D~78_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[23]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[23] .is_wysiwyg = "true";
defparam \instruction_D[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N18
cycloneive_lcell_comb \instruction_EX~8 (
// Equation(s):
// \instruction_EX~8_combout  = (instruction_D[23] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(instruction_D[23]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\branch_taken~0_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\instruction_EX~8_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_EX~8 .lut_mask = 16'h8008;
defparam \instruction_EX~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N13
dffeas \instruction_D[25] (
	.clk(CLK),
	.d(\instruction_D~79_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[25]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[25] .is_wysiwyg = "true";
defparam \instruction_D[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N24
cycloneive_lcell_comb \instruction_EX~9 (
// Equation(s):
// \instruction_EX~9_combout  = (instruction_D[25] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(instruction_D[25]),
	.datab(\branch_taken~0_combout ),
	.datac(\branch_or_jump~2_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\instruction_EX~9_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_EX~9 .lut_mask = 16'h8020;
defparam \instruction_EX~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N6
cycloneive_lcell_comb \ALUOp_EX~0 (
// Equation(s):
// \ALUOp_EX~0_combout  = (\ShiftOp_EX~0_combout  & ((instruction_D[1]) # ((instruction_D[5] & WideOr2)))) # (!\ShiftOp_EX~0_combout  & (instruction_D[5] & ((WideOr2))))

	.dataa(\ShiftOp_EX~0_combout ),
	.datab(instruction_D[5]),
	.datac(instruction_D[1]),
	.datad(\CONTROL_UNIT|WideOr2~0_combout ),
	.cin(gnd),
	.combout(\ALUOp_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~0 .lut_mask = 16'hECA0;
defparam \ALUOp_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N10
cycloneive_lcell_comb \ALUOp_EX~1 (
// Equation(s):
// \ALUOp_EX~1_combout  = (\ALUOp_EX~0_combout  & (!instruction_D[4] & Equal31))

	.dataa(gnd),
	.datab(\ALUOp_EX~0_combout ),
	.datac(instruction_D[4]),
	.datad(\CONTROL_UNIT|Equal3~2_combout ),
	.cin(gnd),
	.combout(\ALUOp_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~1 .lut_mask = 16'h0C00;
defparam \ALUOp_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N10
cycloneive_lcell_comb \ALUOp_EX~2 (
// Equation(s):
// \ALUOp_EX~2_combout  = (!instruction_D[30] & (!instruction_D[31] & !Equal31))

	.dataa(instruction_D[30]),
	.datab(gnd),
	.datac(instruction_D[31]),
	.datad(\CONTROL_UNIT|Equal3~2_combout ),
	.cin(gnd),
	.combout(\ALUOp_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~2 .lut_mask = 16'h0005;
defparam \ALUOp_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N12
cycloneive_lcell_comb \ALUOp_EX~3 (
// Equation(s):
// \ALUOp_EX~3_combout  = (\branch_or_jump~1_combout  & ((\ALUOp_EX~1_combout ) # ((WideOr7 & \ALUOp_EX~2_combout ))))

	.dataa(\ALUOp_EX~1_combout ),
	.datab(\CONTROL_UNIT|WideOr7~0_combout ),
	.datac(\branch_or_jump~1_combout ),
	.datad(\ALUOp_EX~2_combout ),
	.cin(gnd),
	.combout(\ALUOp_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~3 .lut_mask = 16'hE0A0;
defparam \ALUOp_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N18
cycloneive_lcell_comb \ALUOp_EX~4 (
// Equation(s):
// \ALUOp_EX~4_combout  = (instruction_D[26] & (instruction_D[27] & (instruction_D[31] & !instruction_D[28])))

	.dataa(instruction_D[26]),
	.datab(instruction_D[27]),
	.datac(instruction_D[31]),
	.datad(instruction_D[28]),
	.cin(gnd),
	.combout(\ALUOp_EX~4_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~4 .lut_mask = 16'h0080;
defparam \ALUOp_EX~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N24
cycloneive_lcell_comb \ALUOp_EX~5 (
// Equation(s):
// \ALUOp_EX~5_combout  = (\ALUOp_EX~4_combout ) # ((!instruction_D[31] & WideOr6))

	.dataa(instruction_D[31]),
	.datab(\ALUOp_EX~4_combout ),
	.datac(gnd),
	.datad(\CONTROL_UNIT|WideOr6~0_combout ),
	.cin(gnd),
	.combout(\ALUOp_EX~5_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~5 .lut_mask = 16'hDDCC;
defparam \ALUOp_EX~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N6
cycloneive_lcell_comb \ALUOp_EX~6 (
// Equation(s):
// \ALUOp_EX~6_combout  = (\branch_or_jump~1_combout  & (((instruction_D[5] & !WideOr1)) # (!Equal31)))

	.dataa(instruction_D[5]),
	.datab(\CONTROL_UNIT|Equal3~2_combout ),
	.datac(\CONTROL_UNIT|WideOr1~0_combout ),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\ALUOp_EX~6_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~6 .lut_mask = 16'h3B00;
defparam \ALUOp_EX~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N18
cycloneive_lcell_comb \ALUOp_EX~7 (
// Equation(s):
// \ALUOp_EX~7_combout  = (\ALUOp_EX~6_combout  & ((Equal31) # ((\ALUOp_EX~5_combout  & !instruction_D[30]))))

	.dataa(\ALUOp_EX~6_combout ),
	.datab(\ALUOp_EX~5_combout ),
	.datac(\CONTROL_UNIT|Equal3~2_combout ),
	.datad(instruction_D[30]),
	.cin(gnd),
	.combout(\ALUOp_EX~7_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~7 .lut_mask = 16'hA0A8;
defparam \ALUOp_EX~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N24
cycloneive_lcell_comb \ALUOp_EX~8 (
// Equation(s):
// \ALUOp_EX~8_combout  = (instruction_D[5] & (!instruction_D[4] & Equal31))

	.dataa(gnd),
	.datab(instruction_D[5]),
	.datac(instruction_D[4]),
	.datad(\CONTROL_UNIT|Equal3~2_combout ),
	.cin(gnd),
	.combout(\ALUOp_EX~8_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~8 .lut_mask = 16'h0C00;
defparam \ALUOp_EX~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N26
cycloneive_lcell_comb \ALUOp_EX~9 (
// Equation(s):
// \ALUOp_EX~9_combout  = (\ALUOp_EX~8_combout  & (!instruction_D[3] & instruction_D[2]))

	.dataa(gnd),
	.datab(\ALUOp_EX~8_combout ),
	.datac(instruction_D[3]),
	.datad(instruction_D[2]),
	.cin(gnd),
	.combout(\ALUOp_EX~9_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~9 .lut_mask = 16'h0C00;
defparam \ALUOp_EX~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N22
cycloneive_lcell_comb \ALUOp_EX~10 (
// Equation(s):
// \ALUOp_EX~10_combout  = (\branch_or_jump~1_combout  & ((\ALUOp_EX~9_combout ) # ((WideOr5 & \ALUOp_EX~2_combout ))))

	.dataa(\ALUOp_EX~9_combout ),
	.datab(\CONTROL_UNIT|WideOr5~0_combout ),
	.datac(\ALUOp_EX~2_combout ),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\ALUOp_EX~10_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~10 .lut_mask = 16'hEA00;
defparam \ALUOp_EX~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N24
cycloneive_lcell_comb \ALUOp_EX~11 (
// Equation(s):
// \ALUOp_EX~11_combout  = (instruction_D[1] & (instruction_D[3] & (\ALUOp_EX~8_combout  & !instruction_D[2])))

	.dataa(instruction_D[1]),
	.datab(instruction_D[3]),
	.datac(\ALUOp_EX~8_combout ),
	.datad(instruction_D[2]),
	.cin(gnd),
	.combout(\ALUOp_EX~11_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~11 .lut_mask = 16'h0080;
defparam \ALUOp_EX~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N28
cycloneive_lcell_comb \ALUOp_EX~12 (
// Equation(s):
// \ALUOp_EX~12_combout  = (!instruction_D[28] & (instruction_D[27] & (!instruction_D[31] & !instruction_D[30])))

	.dataa(instruction_D[28]),
	.datab(instruction_D[27]),
	.datac(instruction_D[31]),
	.datad(instruction_D[30]),
	.cin(gnd),
	.combout(\ALUOp_EX~12_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~12 .lut_mask = 16'h0004;
defparam \ALUOp_EX~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N12
cycloneive_lcell_comb \ALUOp_EX~13 (
// Equation(s):
// \ALUOp_EX~13_combout  = (\branch_or_jump~1_combout  & ((\ALUOp_EX~11_combout ) # ((\ALUOp_EX~12_combout  & instruction_D[29]))))

	.dataa(\branch_or_jump~1_combout ),
	.datab(\ALUOp_EX~12_combout ),
	.datac(instruction_D[29]),
	.datad(\ALUOp_EX~11_combout ),
	.cin(gnd),
	.combout(\ALUOp_EX~13_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOp_EX~13 .lut_mask = 16'hAA80;
defparam \ALUOp_EX~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N8
cycloneive_lcell_comb \ExtOp_EX~0 (
// Equation(s):
// \ExtOp_EX~0_combout  = (!instruction_D[30] & (!Equal31 & \branch_or_jump~1_combout ))

	.dataa(instruction_D[30]),
	.datab(\CONTROL_UNIT|Equal3~2_combout ),
	.datac(gnd),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\ExtOp_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \ExtOp_EX~0 .lut_mask = 16'h1100;
defparam \ExtOp_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N15
dffeas RegWrite_EX(
	.clk(CLK),
	.d(\RegWrite_EX~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\RegWrite_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam RegWrite_EX.is_wysiwyg = "true";
defparam RegWrite_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N24
cycloneive_lcell_comb \beq_EX~0 (
// Equation(s):
// \beq_EX~0_combout  = (!instruction_D[26] & (!instruction_D[27] & (instruction_D[28] & \j_EX~3_combout )))

	.dataa(instruction_D[26]),
	.datab(instruction_D[27]),
	.datac(instruction_D[28]),
	.datad(\j_EX~3_combout ),
	.cin(gnd),
	.combout(\beq_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \beq_EX~0 .lut_mask = 16'h1000;
defparam \beq_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N30
cycloneive_lcell_comb \bne_EX~0 (
// Equation(s):
// \bne_EX~0_combout  = (instruction_D[26] & (!instruction_D[27] & (instruction_D[28] & \j_EX~3_combout )))

	.dataa(instruction_D[26]),
	.datab(instruction_D[27]),
	.datac(instruction_D[28]),
	.datad(\j_EX~3_combout ),
	.cin(gnd),
	.combout(\bne_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \bne_EX~0 .lut_mask = 16'h2000;
defparam \bne_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N30
cycloneive_lcell_comb \ALUSrc_EX~1 (
// Equation(s):
// \ALUSrc_EX~1_combout  = (\ExtOp_EX~0_combout  & ((instruction_D[29] & ((!WideOr4))) # (!instruction_D[29] & (\ALUOp_EX~4_combout ))))

	.dataa(instruction_D[29]),
	.datab(\ExtOp_EX~0_combout ),
	.datac(\ALUOp_EX~4_combout ),
	.datad(\CONTROL_UNIT|WideOr4~0_combout ),
	.cin(gnd),
	.combout(\ALUSrc_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc_EX~1 .lut_mask = 16'h40C8;
defparam \ALUSrc_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N21
dffeas lui_EX(
	.clk(CLK),
	.d(\lui_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\lui_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam lui_EX.is_wysiwyg = "true";
defparam lui_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N16
cycloneive_lcell_comb \rdata2_EX~8 (
// Equation(s):
// \rdata2_EX~8_combout  = (instruction_D[20] & ((Mux36))) # (!instruction_D[20] & (Mux361))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux36~19_combout ),
	.datad(\REGISTER_FILE|Mux36~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~8 .lut_mask = 16'hFA50;
defparam \rdata2_EX~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N30
cycloneive_lcell_comb \rdata2_EX~9 (
// Equation(s):
// \rdata2_EX~9_combout  = (\always2~2_combout  & ((\rdata2_EX~8_combout ))) # (!\always2~2_combout  & (\portB~29_combout ))

	.dataa(gnd),
	.datab(\portB~29_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~8_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~9_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~9 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N4
cycloneive_lcell_comb \rdata2_EX~12 (
// Equation(s):
// \rdata2_EX~12_combout  = (instruction_D[20] & (Mux38)) # (!instruction_D[20] & ((Mux381)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux38~9_combout ),
	.datad(\REGISTER_FILE|Mux38~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~12 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N20
cycloneive_lcell_comb \rdata2_EX~13 (
// Equation(s):
// \rdata2_EX~13_combout  = (\always2~2_combout  & ((\rdata2_EX~12_combout ))) # (!\always2~2_combout  & (\portB~35_combout ))

	.dataa(\portB~35_combout ),
	.datab(\always2~2_combout ),
	.datac(\rdata2_EX~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdata2_EX~13_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~13 .lut_mask = 16'hE2E2;
defparam \rdata2_EX~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N28
cycloneive_lcell_comb \rdata2_EX~22 (
// Equation(s):
// \rdata2_EX~22_combout  = (instruction_D[20] & (Mux43)) # (!instruction_D[20] & ((Mux431)))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux43~9_combout ),
	.datad(\REGISTER_FILE|Mux43~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~22 .lut_mask = 16'hF3C0;
defparam \rdata2_EX~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N0
cycloneive_lcell_comb \rdata2_EX~23 (
// Equation(s):
// \rdata2_EX~23_combout  = (\always2~2_combout  & ((\rdata2_EX~22_combout ))) # (!\always2~2_combout  & (\portB~50_combout ))

	.dataa(\portB~50_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~22_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~23_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~23 .lut_mask = 16'hFA0A;
defparam \rdata2_EX~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N16
cycloneive_lcell_comb \rdata2_EX~36 (
// Equation(s):
// \rdata2_EX~36_combout  = (instruction_D[20] & (Mux50)) # (!instruction_D[20] & ((Mux501)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux50~9_combout ),
	.datad(\REGISTER_FILE|Mux50~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~36_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~36 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N28
cycloneive_lcell_comb \rdata2_EX~37 (
// Equation(s):
// \rdata2_EX~37_combout  = (\always2~2_combout  & ((\rdata2_EX~36_combout ))) # (!\always2~2_combout  & (\portB~68_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portB~68_combout ),
	.datad(\rdata2_EX~36_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~37_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~37 .lut_mask = 16'hFC30;
defparam \rdata2_EX~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N18
cycloneive_lcell_comb \rdata2_EX~42 (
// Equation(s):
// \rdata2_EX~42_combout  = (instruction_D[20] & (Mux55)) # (!instruction_D[20] & ((Mux551)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux55~9_combout ),
	.datad(\REGISTER_FILE|Mux55~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~42_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~42 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N4
cycloneive_lcell_comb \rdata2_EX~43 (
// Equation(s):
// \rdata2_EX~43_combout  = (\always2~2_combout  & ((\rdata2_EX~42_combout ))) # (!\always2~2_combout  & (\portB~76_combout ))

	.dataa(gnd),
	.datab(\portB~76_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~42_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~43_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~43 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N5
dffeas \instruction_D[11] (
	.clk(CLK),
	.d(\instruction_D~92_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[11]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[11] .is_wysiwyg = "true";
defparam \instruction_D[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N28
cycloneive_lcell_comb \imm_EX~6 (
// Equation(s):
// \imm_EX~6_combout  = (instruction_D[11] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(instruction_D[11]),
	.datac(\branch_taken~0_combout ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\imm_EX~6_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~6 .lut_mask = 16'h8400;
defparam \imm_EX~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N2
cycloneive_lcell_comb \rdata2_EX~44 (
// Equation(s):
// \rdata2_EX~44_combout  = (instruction_D[20] & ((Mux52))) # (!instruction_D[20] & (Mux521))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux52~19_combout ),
	.datad(\REGISTER_FILE|Mux52~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~44_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~44 .lut_mask = 16'hFC30;
defparam \rdata2_EX~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N26
cycloneive_lcell_comb \rdata2_EX~45 (
// Equation(s):
// \rdata2_EX~45_combout  = (\always2~2_combout  & ((\rdata2_EX~44_combout ))) # (!\always2~2_combout  & (\portB~108_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portB~108_combout ),
	.datad(\rdata2_EX~44_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~45_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~45 .lut_mask = 16'hFC30;
defparam \rdata2_EX~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N30
cycloneive_lcell_comb \rdata2_EX~46 (
// Equation(s):
// \rdata2_EX~46_combout  = (instruction_D[20] & (Mux53)) # (!instruction_D[20] & ((Mux531)))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux53~9_combout ),
	.datad(\REGISTER_FILE|Mux53~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~46_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~46 .lut_mask = 16'hF3C0;
defparam \rdata2_EX~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N18
cycloneive_lcell_comb \rdata2_EX~47 (
// Equation(s):
// \rdata2_EX~47_combout  = (\always2~2_combout  & ((\rdata2_EX~46_combout ))) # (!\always2~2_combout  & (\portB~109_combout ))

	.dataa(\portB~109_combout ),
	.datab(\always2~2_combout ),
	.datac(\rdata2_EX~46_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdata2_EX~47_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~47 .lut_mask = 16'hE2E2;
defparam \rdata2_EX~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N10
cycloneive_lcell_comb \rdata2_EX~48 (
// Equation(s):
// \rdata2_EX~48_combout  = (instruction_D[20] & ((Mux56))) # (!instruction_D[20] & (Mux561))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux56~19_combout ),
	.datad(\REGISTER_FILE|Mux56~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~48_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~48 .lut_mask = 16'hFC30;
defparam \rdata2_EX~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N28
cycloneive_lcell_comb \rdata2_EX~49 (
// Equation(s):
// \rdata2_EX~49_combout  = (\always2~2_combout  & ((\rdata2_EX~48_combout ))) # (!\always2~2_combout  & (\portB~82_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portB~82_combout ),
	.datad(\rdata2_EX~48_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~49_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~49 .lut_mask = 16'hFC30;
defparam \rdata2_EX~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N2
cycloneive_lcell_comb \rdata2_EX~52 (
// Equation(s):
// \rdata2_EX~52_combout  = (instruction_D[20] & ((Mux58))) # (!instruction_D[20] & (Mux581))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux58~19_combout ),
	.datad(\REGISTER_FILE|Mux58~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~52_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~52 .lut_mask = 16'hFC30;
defparam \rdata2_EX~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N28
cycloneive_lcell_comb \rdata2_EX~53 (
// Equation(s):
// \rdata2_EX~53_combout  = (\always2~2_combout  & ((\rdata2_EX~52_combout ))) # (!\always2~2_combout  & (\portB~87_combout ))

	.dataa(gnd),
	.datab(\portB~87_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~52_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~53_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~53 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N22
cycloneive_lcell_comb \rdata1_EX~2 (
// Equation(s):
// \rdata1_EX~2_combout  = (instruction_D[25] & (Mux29)) # (!instruction_D[25] & ((Mux291)))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux29~9_combout ),
	.datad(\REGISTER_FILE|Mux29~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~2 .lut_mask = 16'hF5A0;
defparam \rdata1_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N4
cycloneive_lcell_comb \rdata1_EX~3 (
// Equation(s):
// \rdata1_EX~3_combout  = (\always2~2_combout  & ((\rdata1_EX~2_combout ))) # (!\always2~2_combout  & (\portA~9_combout ))

	.dataa(gnd),
	.datab(\portA~9_combout ),
	.datac(\rdata1_EX~2_combout ),
	.datad(\always2~2_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~3 .lut_mask = 16'hF0CC;
defparam \rdata1_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N6
cycloneive_lcell_comb \rdata1_EX~4 (
// Equation(s):
// \rdata1_EX~4_combout  = (instruction_D[25] & (Mux30)) # (!instruction_D[25] & ((Mux301)))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux30~9_combout ),
	.datad(\REGISTER_FILE|Mux30~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~4 .lut_mask = 16'hF5A0;
defparam \rdata1_EX~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N10
cycloneive_lcell_comb \rdata1_EX~5 (
// Equation(s):
// \rdata1_EX~5_combout  = (\always2~2_combout  & ((\rdata1_EX~4_combout ))) # (!\always2~2_combout  & (\portA~12_combout ))

	.dataa(\portA~12_combout ),
	.datab(\always2~2_combout ),
	.datac(\rdata1_EX~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdata1_EX~5_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~5 .lut_mask = 16'hE2E2;
defparam \rdata1_EX~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N20
cycloneive_lcell_comb \rdata2_EX~54 (
// Equation(s):
// \rdata2_EX~54_combout  = (instruction_D[20] & (Mux63)) # (!instruction_D[20] & ((Mux631)))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux63~9_combout ),
	.datad(\REGISTER_FILE|Mux63~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~54_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~54 .lut_mask = 16'hF3C0;
defparam \rdata2_EX~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N6
cycloneive_lcell_comb \rdata2_EX~55 (
// Equation(s):
// \rdata2_EX~55_combout  = (\always2~2_combout  & ((\rdata2_EX~54_combout ))) # (!\always2~2_combout  & (\portB~92_combout ))

	.dataa(\portB~92_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata2_EX~54_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~55_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~55 .lut_mask = 16'hEE22;
defparam \rdata2_EX~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N18
cycloneive_lcell_comb \rdata2_EX~56 (
// Equation(s):
// \rdata2_EX~56_combout  = (instruction_D[20] & (Mux62)) # (!instruction_D[20] & ((Mux621)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux62~9_combout ),
	.datad(\REGISTER_FILE|Mux62~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~56_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~56 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N0
cycloneive_lcell_comb \rdata2_EX~57 (
// Equation(s):
// \rdata2_EX~57_combout  = (\always2~2_combout  & ((\rdata2_EX~56_combout ))) # (!\always2~2_combout  & (\portB~97_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portB~97_combout ),
	.datad(\rdata2_EX~56_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~57_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~57 .lut_mask = 16'hFC30;
defparam \rdata2_EX~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N0
cycloneive_lcell_comb \rdata1_EX~6 (
// Equation(s):
// \rdata1_EX~6_combout  = (instruction_D[25] & ((Mux27))) # (!instruction_D[25] & (Mux271))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux27~19_combout ),
	.datad(\REGISTER_FILE|Mux27~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~6 .lut_mask = 16'hFC30;
defparam \rdata1_EX~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N24
cycloneive_lcell_comb \rdata1_EX~7 (
// Equation(s):
// \rdata1_EX~7_combout  = (\always2~2_combout  & ((\rdata1_EX~6_combout ))) # (!\always2~2_combout  & (\portA~14_combout ))

	.dataa(gnd),
	.datab(\portA~14_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~6_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~7_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~7 .lut_mask = 16'hFC0C;
defparam \rdata1_EX~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N6
cycloneive_lcell_comb \rdata1_EX~8 (
// Equation(s):
// \rdata1_EX~8_combout  = (instruction_D[25] & (Mux28)) # (!instruction_D[25] & ((Mux281)))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux28~9_combout ),
	.datad(\REGISTER_FILE|Mux28~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~8 .lut_mask = 16'hF5A0;
defparam \rdata1_EX~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N28
cycloneive_lcell_comb \rdata1_EX~9 (
// Equation(s):
// \rdata1_EX~9_combout  = (\always2~2_combout  & ((\rdata1_EX~8_combout ))) # (!\always2~2_combout  & (\portA~16_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portA~16_combout ),
	.datad(\rdata1_EX~8_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~9_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~9 .lut_mask = 16'hFC30;
defparam \rdata1_EX~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N0
cycloneive_lcell_comb \rdata1_EX~10 (
// Equation(s):
// \rdata1_EX~10_combout  = (instruction_D[25] & ((Mux23))) # (!instruction_D[25] & (Mux231))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux23~19_combout ),
	.datad(\REGISTER_FILE|Mux23~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~10 .lut_mask = 16'hFA50;
defparam \rdata1_EX~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N14
cycloneive_lcell_comb \rdata1_EX~11 (
// Equation(s):
// \rdata1_EX~11_combout  = (\always2~2_combout  & ((\rdata1_EX~10_combout ))) # (!\always2~2_combout  & (\portA~17_combout ))

	.dataa(gnd),
	.datab(\portA~17_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~10_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~11_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~11 .lut_mask = 16'hFC0C;
defparam \rdata1_EX~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N22
cycloneive_lcell_comb \rdata1_EX~12 (
// Equation(s):
// \rdata1_EX~12_combout  = (instruction_D[25] & ((Mux24))) # (!instruction_D[25] & (Mux241))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux24~19_combout ),
	.datad(\REGISTER_FILE|Mux24~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~12 .lut_mask = 16'hFA50;
defparam \rdata1_EX~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N0
cycloneive_lcell_comb \rdata1_EX~13 (
// Equation(s):
// \rdata1_EX~13_combout  = (\always2~2_combout  & ((\rdata1_EX~12_combout ))) # (!\always2~2_combout  & (\portA~19_combout ))

	.dataa(\portA~19_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata1_EX~12_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~13_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~13 .lut_mask = 16'hEE22;
defparam \rdata1_EX~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N28
cycloneive_lcell_comb \rdata1_EX~14 (
// Equation(s):
// \rdata1_EX~14_combout  = (instruction_D[25] & (Mux25)) # (!instruction_D[25] & ((Mux251)))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux25~9_combout ),
	.datad(\REGISTER_FILE|Mux25~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~14 .lut_mask = 16'hF3C0;
defparam \rdata1_EX~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N2
cycloneive_lcell_comb \rdata1_EX~15 (
// Equation(s):
// \rdata1_EX~15_combout  = (\always2~2_combout  & ((\rdata1_EX~14_combout ))) # (!\always2~2_combout  & (\portA~21_combout ))

	.dataa(\portA~21_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata1_EX~14_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~15_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~15 .lut_mask = 16'hEE22;
defparam \rdata1_EX~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N16
cycloneive_lcell_comb \rdata1_EX~16 (
// Equation(s):
// \rdata1_EX~16_combout  = (instruction_D[25] & ((Mux26))) # (!instruction_D[25] & (Mux261))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux26~19_combout ),
	.datad(\REGISTER_FILE|Mux26~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~16 .lut_mask = 16'hFC30;
defparam \rdata1_EX~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N8
cycloneive_lcell_comb \rdata1_EX~17 (
// Equation(s):
// \rdata1_EX~17_combout  = (\always2~2_combout  & ((\rdata1_EX~16_combout ))) # (!\always2~2_combout  & (\portA~23_combout ))

	.dataa(\portA~23_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata1_EX~16_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~17_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~17 .lut_mask = 16'hEE22;
defparam \rdata1_EX~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N2
cycloneive_lcell_comb \rdata2_EX~60 (
// Equation(s):
// \rdata2_EX~60_combout  = (instruction_D[20] & (Mux60)) # (!instruction_D[20] & ((Mux601)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux60~9_combout ),
	.datad(\REGISTER_FILE|Mux60~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~60_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~60 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N30
cycloneive_lcell_comb \rdata2_EX~61 (
// Equation(s):
// \rdata2_EX~61_combout  = (\always2~2_combout  & ((\rdata2_EX~60_combout ))) # (!\always2~2_combout  & (\portB~103_combout ))

	.dataa(\portB~103_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~60_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~61_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~61 .lut_mask = 16'hFA0A;
defparam \rdata2_EX~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N0
cycloneive_lcell_comb \rdata1_EX~18 (
// Equation(s):
// \rdata1_EX~18_combout  = (instruction_D[25] & ((Mux15))) # (!instruction_D[25] & (Mux151))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux15~19_combout ),
	.datad(\REGISTER_FILE|Mux15~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~18 .lut_mask = 16'hFC30;
defparam \rdata1_EX~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N30
cycloneive_lcell_comb \rdata1_EX~19 (
// Equation(s):
// \rdata1_EX~19_combout  = (\always2~2_combout  & ((\rdata1_EX~18_combout ))) # (!\always2~2_combout  & (\portA~25_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portA~25_combout ),
	.datad(\rdata1_EX~18_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~19_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~19 .lut_mask = 16'hFC30;
defparam \rdata1_EX~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N10
cycloneive_lcell_comb \rdata1_EX~20 (
// Equation(s):
// \rdata1_EX~20_combout  = (instruction_D[25] & (Mux16)) # (!instruction_D[25] & ((Mux161)))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux16~9_combout ),
	.datad(\REGISTER_FILE|Mux16~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~20 .lut_mask = 16'hF3C0;
defparam \rdata1_EX~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N4
cycloneive_lcell_comb \rdata1_EX~21 (
// Equation(s):
// \rdata1_EX~21_combout  = (\always2~2_combout  & ((\rdata1_EX~20_combout ))) # (!\always2~2_combout  & (\portA~27_combout ))

	.dataa(\portA~27_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata1_EX~20_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~21_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~21 .lut_mask = 16'hEE22;
defparam \rdata1_EX~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N10
cycloneive_lcell_comb \rdata1_EX~22 (
// Equation(s):
// \rdata1_EX~22_combout  = (instruction_D[25] & ((Mux17))) # (!instruction_D[25] & (Mux171))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux17~19_combout ),
	.datad(\REGISTER_FILE|Mux17~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~22 .lut_mask = 16'hFA50;
defparam \rdata1_EX~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N4
cycloneive_lcell_comb \rdata1_EX~23 (
// Equation(s):
// \rdata1_EX~23_combout  = (\always2~2_combout  & ((\rdata1_EX~22_combout ))) # (!\always2~2_combout  & (\portA~29_combout ))

	.dataa(gnd),
	.datab(\portA~29_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~22_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~23_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~23 .lut_mask = 16'hFC0C;
defparam \rdata1_EX~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N20
cycloneive_lcell_comb \rdata1_EX~24 (
// Equation(s):
// \rdata1_EX~24_combout  = (instruction_D[25] & (Mux18)) # (!instruction_D[25] & ((Mux181)))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux18~9_combout ),
	.datad(\REGISTER_FILE|Mux18~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~24 .lut_mask = 16'hF5A0;
defparam \rdata1_EX~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N18
cycloneive_lcell_comb \rdata1_EX~25 (
// Equation(s):
// \rdata1_EX~25_combout  = (\always2~2_combout  & ((\rdata1_EX~24_combout ))) # (!\always2~2_combout  & (\portA~31_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portA~31_combout ),
	.datad(\rdata1_EX~24_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~25_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~25 .lut_mask = 16'hFC30;
defparam \rdata1_EX~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N12
cycloneive_lcell_comb \rdata1_EX~26 (
// Equation(s):
// \rdata1_EX~26_combout  = (instruction_D[25] & ((Mux19))) # (!instruction_D[25] & (Mux191))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux19~19_combout ),
	.datad(\REGISTER_FILE|Mux19~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~26 .lut_mask = 16'hFA50;
defparam \rdata1_EX~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N8
cycloneive_lcell_comb \rdata1_EX~27 (
// Equation(s):
// \rdata1_EX~27_combout  = (\always2~2_combout  & ((\rdata1_EX~26_combout ))) # (!\always2~2_combout  & (\portA~33_combout ))

	.dataa(gnd),
	.datab(\portA~33_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~26_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~27_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~27 .lut_mask = 16'hFC0C;
defparam \rdata1_EX~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N22
cycloneive_lcell_comb \rdata1_EX~28 (
// Equation(s):
// \rdata1_EX~28_combout  = (instruction_D[25] & ((Mux20))) # (!instruction_D[25] & (Mux201))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux20~19_combout ),
	.datad(\REGISTER_FILE|Mux20~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~28 .lut_mask = 16'hFC30;
defparam \rdata1_EX~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N6
cycloneive_lcell_comb \rdata1_EX~29 (
// Equation(s):
// \rdata1_EX~29_combout  = (\always2~2_combout  & ((\rdata1_EX~28_combout ))) # (!\always2~2_combout  & (\portA~35_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portA~35_combout ),
	.datad(\rdata1_EX~28_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~29_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~29 .lut_mask = 16'hFC30;
defparam \rdata1_EX~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N18
cycloneive_lcell_comb \rdata1_EX~30 (
// Equation(s):
// \rdata1_EX~30_combout  = (instruction_D[25] & ((Mux21))) # (!instruction_D[25] & (Mux211))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux21~19_combout ),
	.datad(\REGISTER_FILE|Mux21~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~30 .lut_mask = 16'hFA50;
defparam \rdata1_EX~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N2
cycloneive_lcell_comb \rdata1_EX~31 (
// Equation(s):
// \rdata1_EX~31_combout  = (\always2~2_combout  & ((\rdata1_EX~30_combout ))) # (!\always2~2_combout  & (\portA~36_combout ))

	.dataa(\portA~36_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~30_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~31_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~31 .lut_mask = 16'hFA0A;
defparam \rdata1_EX~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N12
cycloneive_lcell_comb \rdata1_EX~32 (
// Equation(s):
// \rdata1_EX~32_combout  = (instruction_D[25] & (Mux22)) # (!instruction_D[25] & ((Mux221)))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux22~9_combout ),
	.datad(\REGISTER_FILE|Mux22~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~32_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~32 .lut_mask = 16'hF5A0;
defparam \rdata1_EX~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N28
cycloneive_lcell_comb \rdata1_EX~33 (
// Equation(s):
// \rdata1_EX~33_combout  = (\always2~2_combout  & ((\rdata1_EX~32_combout ))) # (!\always2~2_combout  & (\portA~37_combout ))

	.dataa(gnd),
	.datab(\portA~37_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~32_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~33_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~33 .lut_mask = 16'hFC0C;
defparam \rdata1_EX~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N22
cycloneive_lcell_comb \rdata1_EX~34 (
// Equation(s):
// \rdata1_EX~34_combout  = (instruction_D[25] & ((Mux0))) # (!instruction_D[25] & (Mux01))

	.dataa(instruction_D[25]),
	.datab(\REGISTER_FILE|Mux0~19_combout ),
	.datac(\REGISTER_FILE|Mux0~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdata1_EX~34_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~34 .lut_mask = 16'hE4E4;
defparam \rdata1_EX~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N14
cycloneive_lcell_comb \rdata1_EX~35 (
// Equation(s):
// \rdata1_EX~35_combout  = (\always2~2_combout  & ((\rdata1_EX~34_combout ))) # (!\always2~2_combout  & (\portA~39_combout ))

	.dataa(\portA~39_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~34_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~35_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~35 .lut_mask = 16'hFA0A;
defparam \rdata1_EX~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N14
cycloneive_lcell_comb \rdata1_EX~36 (
// Equation(s):
// \rdata1_EX~36_combout  = (instruction_D[25] & ((Mux2))) # (!instruction_D[25] & (Mux210))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux2~19_combout ),
	.datad(\REGISTER_FILE|Mux2~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~36_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~36 .lut_mask = 16'hFA50;
defparam \rdata1_EX~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N24
cycloneive_lcell_comb \rdata1_EX~37 (
// Equation(s):
// \rdata1_EX~37_combout  = (\always2~2_combout  & ((\rdata1_EX~36_combout ))) # (!\always2~2_combout  & (\portA~41_combout ))

	.dataa(gnd),
	.datab(\portA~41_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~36_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~37_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~37 .lut_mask = 16'hFC0C;
defparam \rdata1_EX~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N30
cycloneive_lcell_comb \rdata1_EX~38 (
// Equation(s):
// \rdata1_EX~38_combout  = (instruction_D[25] & ((Mux1))) # (!instruction_D[25] & (Mux11))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux1~19_combout ),
	.datad(\REGISTER_FILE|Mux1~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~38_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~38 .lut_mask = 16'hFA50;
defparam \rdata1_EX~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N22
cycloneive_lcell_comb \rdata1_EX~39 (
// Equation(s):
// \rdata1_EX~39_combout  = (\always2~2_combout  & ((\rdata1_EX~38_combout ))) # (!\always2~2_combout  & (\portA~43_combout ))

	.dataa(\portA~43_combout ),
	.datab(\always2~2_combout ),
	.datac(\rdata1_EX~38_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdata1_EX~39_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~39 .lut_mask = 16'hE2E2;
defparam \rdata1_EX~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N30
cycloneive_lcell_comb \rdata1_EX~40 (
// Equation(s):
// \rdata1_EX~40_combout  = (instruction_D[25] & (Mux3)) # (!instruction_D[25] & ((Mux31)))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux3~9_combout ),
	.datad(\REGISTER_FILE|Mux3~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~40_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~40 .lut_mask = 16'hF5A0;
defparam \rdata1_EX~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N28
cycloneive_lcell_comb \rdata1_EX~41 (
// Equation(s):
// \rdata1_EX~41_combout  = (\always2~2_combout  & ((\rdata1_EX~40_combout ))) # (!\always2~2_combout  & (\portA~45_combout ))

	.dataa(gnd),
	.datab(\portA~45_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~40_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~41_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~41 .lut_mask = 16'hFC0C;
defparam \rdata1_EX~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N0
cycloneive_lcell_comb \rdata1_EX~42 (
// Equation(s):
// \rdata1_EX~42_combout  = (instruction_D[25] & (Mux4)) # (!instruction_D[25] & ((Mux410)))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux4~9_combout ),
	.datad(\REGISTER_FILE|Mux4~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~42_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~42 .lut_mask = 16'hF3C0;
defparam \rdata1_EX~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N4
cycloneive_lcell_comb \rdata1_EX~43 (
// Equation(s):
// \rdata1_EX~43_combout  = (\always2~2_combout  & ((\rdata1_EX~42_combout ))) # (!\always2~2_combout  & (\portA~47_combout ))

	.dataa(\portA~47_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata1_EX~42_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~43_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~43 .lut_mask = 16'hEE22;
defparam \rdata1_EX~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N10
cycloneive_lcell_comb \rdata1_EX~44 (
// Equation(s):
// \rdata1_EX~44_combout  = (instruction_D[25] & ((Mux5))) # (!instruction_D[25] & (Mux510))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux5~19_combout ),
	.datad(\REGISTER_FILE|Mux5~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~44_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~44 .lut_mask = 16'hFA50;
defparam \rdata1_EX~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N20
cycloneive_lcell_comb \rdata1_EX~45 (
// Equation(s):
// \rdata1_EX~45_combout  = (\always2~2_combout  & ((\rdata1_EX~44_combout ))) # (!\always2~2_combout  & (\portA~49_combout ))

	.dataa(\portA~49_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~44_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~45_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~45 .lut_mask = 16'hFA0A;
defparam \rdata1_EX~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N30
cycloneive_lcell_comb \rdata1_EX~46 (
// Equation(s):
// \rdata1_EX~46_combout  = (instruction_D[25] & (Mux6)) # (!instruction_D[25] & ((Mux64)))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux6~9_combout ),
	.datad(\REGISTER_FILE|Mux6~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~46_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~46 .lut_mask = 16'hF3C0;
defparam \rdata1_EX~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N6
cycloneive_lcell_comb \rdata1_EX~47 (
// Equation(s):
// \rdata1_EX~47_combout  = (\always2~2_combout  & ((\rdata1_EX~46_combout ))) # (!\always2~2_combout  & (\portA~51_combout ))

	.dataa(gnd),
	.datab(\portA~51_combout ),
	.datac(\rdata1_EX~46_combout ),
	.datad(\always2~2_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~47_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~47 .lut_mask = 16'hF0CC;
defparam \rdata1_EX~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N30
cycloneive_lcell_comb \rdata1_EX~48 (
// Equation(s):
// \rdata1_EX~48_combout  = (instruction_D[25] & ((Mux7))) # (!instruction_D[25] & (Mux71))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux7~19_combout ),
	.datad(\REGISTER_FILE|Mux7~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~48_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~48 .lut_mask = 16'hFA50;
defparam \rdata1_EX~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N30
cycloneive_lcell_comb \rdata1_EX~49 (
// Equation(s):
// \rdata1_EX~49_combout  = (\always2~2_combout  & ((\rdata1_EX~48_combout ))) # (!\always2~2_combout  & (\portA~53_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portA~53_combout ),
	.datad(\rdata1_EX~48_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~49_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~49 .lut_mask = 16'hFC30;
defparam \rdata1_EX~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N12
cycloneive_lcell_comb \rdata1_EX~50 (
// Equation(s):
// \rdata1_EX~50_combout  = (instruction_D[25] & (Mux8)) # (!instruction_D[25] & ((Mux81)))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux8~9_combout ),
	.datad(\REGISTER_FILE|Mux8~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~50_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~50 .lut_mask = 16'hF3C0;
defparam \rdata1_EX~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N20
cycloneive_lcell_comb \rdata1_EX~51 (
// Equation(s):
// \rdata1_EX~51_combout  = (\always2~2_combout  & ((\rdata1_EX~50_combout ))) # (!\always2~2_combout  & (\portA~55_combout ))

	.dataa(\portA~55_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata1_EX~50_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~51_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~51 .lut_mask = 16'hEE22;
defparam \rdata1_EX~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N14
cycloneive_lcell_comb \rdata1_EX~52 (
// Equation(s):
// \rdata1_EX~52_combout  = (instruction_D[25] & (Mux9)) # (!instruction_D[25] & ((Mux91)))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux9~9_combout ),
	.datad(\REGISTER_FILE|Mux9~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~52_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~52 .lut_mask = 16'hF3C0;
defparam \rdata1_EX~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N8
cycloneive_lcell_comb \rdata1_EX~53 (
// Equation(s):
// \rdata1_EX~53_combout  = (\always2~2_combout  & ((\rdata1_EX~52_combout ))) # (!\always2~2_combout  & (\portA~57_combout ))

	.dataa(\portA~57_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~52_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~53_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~53 .lut_mask = 16'hFA0A;
defparam \rdata1_EX~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N20
cycloneive_lcell_comb \rdata1_EX~54 (
// Equation(s):
// \rdata1_EX~54_combout  = (instruction_D[25] & ((Mux10))) # (!instruction_D[25] & (Mux101))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux10~19_combout ),
	.datad(\REGISTER_FILE|Mux10~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~54_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~54 .lut_mask = 16'hFC30;
defparam \rdata1_EX~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N30
cycloneive_lcell_comb \rdata1_EX~55 (
// Equation(s):
// \rdata1_EX~55_combout  = (\always2~2_combout  & ((\rdata1_EX~54_combout ))) # (!\always2~2_combout  & (\portA~59_combout ))

	.dataa(\portA~59_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata1_EX~54_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~55_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~55 .lut_mask = 16'hEE22;
defparam \rdata1_EX~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N16
cycloneive_lcell_comb \rdata1_EX~56 (
// Equation(s):
// \rdata1_EX~56_combout  = (instruction_D[25] & (Mux111)) # (!instruction_D[25] & ((Mux112)))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux11~9_combout ),
	.datad(\REGISTER_FILE|Mux11~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~56_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~56 .lut_mask = 16'hF5A0;
defparam \rdata1_EX~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N26
cycloneive_lcell_comb \rdata1_EX~57 (
// Equation(s):
// \rdata1_EX~57_combout  = (\always2~2_combout  & ((\rdata1_EX~56_combout ))) # (!\always2~2_combout  & (\portA~61_combout ))

	.dataa(gnd),
	.datab(\portA~61_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~56_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~57_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~57 .lut_mask = 16'hFC0C;
defparam \rdata1_EX~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N14
cycloneive_lcell_comb \rdata1_EX~58 (
// Equation(s):
// \rdata1_EX~58_combout  = (instruction_D[25] & (Mux12)) # (!instruction_D[25] & ((Mux121)))

	.dataa(gnd),
	.datab(instruction_D[25]),
	.datac(\REGISTER_FILE|Mux12~9_combout ),
	.datad(\REGISTER_FILE|Mux12~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~58_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~58 .lut_mask = 16'hF3C0;
defparam \rdata1_EX~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N18
cycloneive_lcell_comb \rdata1_EX~59 (
// Equation(s):
// \rdata1_EX~59_combout  = (\always2~2_combout  & ((\rdata1_EX~58_combout ))) # (!\always2~2_combout  & (\portA~63_combout ))

	.dataa(\portA~63_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata1_EX~58_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~59_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~59 .lut_mask = 16'hFA0A;
defparam \rdata1_EX~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N28
cycloneive_lcell_comb \rdata1_EX~60 (
// Equation(s):
// \rdata1_EX~60_combout  = (instruction_D[25] & (Mux13)) # (!instruction_D[25] & ((Mux131)))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux13~9_combout ),
	.datad(\REGISTER_FILE|Mux13~19_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~60_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~60 .lut_mask = 16'hF5A0;
defparam \rdata1_EX~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N2
cycloneive_lcell_comb \rdata1_EX~61 (
// Equation(s):
// \rdata1_EX~61_combout  = (\always2~2_combout  & ((\rdata1_EX~60_combout ))) # (!\always2~2_combout  & (\portA~65_combout ))

	.dataa(\portA~65_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata1_EX~60_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~61_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~61 .lut_mask = 16'hEE22;
defparam \rdata1_EX~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N18
cycloneive_lcell_comb \rdata1_EX~62 (
// Equation(s):
// \rdata1_EX~62_combout  = (instruction_D[25] & ((Mux14))) # (!instruction_D[25] & (Mux141))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux14~19_combout ),
	.datad(\REGISTER_FILE|Mux14~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~62_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~62 .lut_mask = 16'hFA50;
defparam \rdata1_EX~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N12
cycloneive_lcell_comb \rdata1_EX~63 (
// Equation(s):
// \rdata1_EX~63_combout  = (\always2~2_combout  & ((\rdata1_EX~62_combout ))) # (!\always2~2_combout  & (\portA~67_combout ))

	.dataa(\portA~67_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata1_EX~62_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~63_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~63 .lut_mask = 16'hEE22;
defparam \rdata1_EX~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N28
cycloneive_lcell_comb \Decoder0~0 (
// Equation(s):
// \Decoder0~0_combout  = (\Add2~2_combout  & !\Add2~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~2_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~0 .lut_mask = 16'h00F0;
defparam \Decoder0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N6
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (\Add2~2_combout  & (((\Add2~0_combout )))) # (!\Add2~2_combout  & ((\Add2~0_combout  & (\btbframes.frameblocks[1].tag [15])) # (!\Add2~0_combout  & ((\btbframes.frameblocks[0].tag [15])))))

	.dataa(\btbframes.frameblocks[1].tag [15]),
	.datab(\Add2~2_combout ),
	.datac(\Add2~0_combout ),
	.datad(\btbframes.frameblocks[0].tag [15]),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hE3E0;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N24
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (\Add2~2_combout  & ((\Mux13~0_combout  & (\btbframes.frameblocks[3].tag [15])) # (!\Mux13~0_combout  & ((\btbframes.frameblocks[2].tag [15]))))) # (!\Add2~2_combout  & (((\Mux13~0_combout ))))

	.dataa(\btbframes.frameblocks[3].tag [15]),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[2].tag [15]),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hBBC0;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N28
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (\Add2~0_combout  & (\Add2~2_combout )) # (!\Add2~0_combout  & ((\Add2~2_combout  & (\btbframes.frameblocks[2].tag [16])) # (!\Add2~2_combout  & ((\btbframes.frameblocks[0].tag [16])))))

	.dataa(\Add2~0_combout ),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[2].tag [16]),
	.datad(\btbframes.frameblocks[0].tag [16]),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hD9C8;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N14
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (\Add2~0_combout  & ((\Mux12~0_combout  & (\btbframes.frameblocks[3].tag [16])) # (!\Mux12~0_combout  & ((\btbframes.frameblocks[1].tag [16]))))) # (!\Add2~0_combout  & (((\Mux12~0_combout ))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[3].tag [16]),
	.datac(\btbframes.frameblocks[1].tag [16]),
	.datad(\Mux12~0_combout ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hDDA0;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N12
cycloneive_lcell_comb \does_exist~0 (
// Equation(s):
// \does_exist~0_combout  = (\Mux13~1_combout  & (\Add2~34_combout  & (\Mux12~1_combout  $ (!\Add2~36_combout )))) # (!\Mux13~1_combout  & (!\Add2~34_combout  & (\Mux12~1_combout  $ (!\Add2~36_combout ))))

	.dataa(\Mux13~1_combout ),
	.datab(\Add2~34_combout ),
	.datac(\Mux12~1_combout ),
	.datad(\Add2~36_combout ),
	.cin(gnd),
	.combout(\does_exist~0_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~0 .lut_mask = 16'h9009;
defparam \does_exist~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N12
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (\Add2~0_combout  & ((\btbframes.frameblocks[1].tag [17]) # ((\Add2~2_combout )))) # (!\Add2~0_combout  & (((!\Add2~2_combout  & \btbframes.frameblocks[0].tag [17]))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[1].tag [17]),
	.datac(\Add2~2_combout ),
	.datad(\btbframes.frameblocks[0].tag [17]),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hADA8;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N18
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (\Add2~2_combout  & ((\Mux11~0_combout  & ((\btbframes.frameblocks[3].tag [17]))) # (!\Mux11~0_combout  & (\btbframes.frameblocks[2].tag [17])))) # (!\Add2~2_combout  & (((\Mux11~0_combout ))))

	.dataa(\btbframes.frameblocks[2].tag [17]),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[3].tag [17]),
	.datad(\Mux11~0_combout ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hF388;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N22
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (\Add2~2_combout  & (((\btbframes.frameblocks[2].tag [18]) # (\Add2~0_combout )))) # (!\Add2~2_combout  & (\btbframes.frameblocks[0].tag [18] & ((!\Add2~0_combout ))))

	.dataa(\btbframes.frameblocks[0].tag [18]),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[2].tag [18]),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hCCE2;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N8
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (\Add2~0_combout  & ((\Mux10~0_combout  & (\btbframes.frameblocks[3].tag [18])) # (!\Mux10~0_combout  & ((\btbframes.frameblocks[1].tag [18]))))) # (!\Add2~0_combout  & (((\Mux10~0_combout ))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[3].tag [18]),
	.datac(\Mux10~0_combout ),
	.datad(\btbframes.frameblocks[1].tag [18]),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hDAD0;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N18
cycloneive_lcell_comb \does_exist~1 (
// Equation(s):
// \does_exist~1_combout  = (\Mux11~1_combout  & (\Add2~38_combout  & (\Add2~40_combout  $ (!\Mux10~1_combout )))) # (!\Mux11~1_combout  & (!\Add2~38_combout  & (\Add2~40_combout  $ (!\Mux10~1_combout ))))

	.dataa(\Mux11~1_combout ),
	.datab(\Add2~40_combout ),
	.datac(\Mux10~1_combout ),
	.datad(\Add2~38_combout ),
	.cin(gnd),
	.combout(\does_exist~1_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~1 .lut_mask = 16'h8241;
defparam \does_exist~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N16
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (\Add2~0_combout  & ((\btbframes.frameblocks[1].tag [19]) # ((\Add2~2_combout )))) # (!\Add2~0_combout  & (((!\Add2~2_combout  & \btbframes.frameblocks[0].tag [19]))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[1].tag [19]),
	.datac(\Add2~2_combout ),
	.datad(\btbframes.frameblocks[0].tag [19]),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hADA8;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N2
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (\Add2~2_combout  & ((\Mux9~0_combout  & ((\btbframes.frameblocks[3].tag [19]))) # (!\Mux9~0_combout  & (\btbframes.frameblocks[2].tag [19])))) # (!\Add2~2_combout  & (((\Mux9~0_combout ))))

	.dataa(\btbframes.frameblocks[2].tag [19]),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[3].tag [19]),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hF388;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N0
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (\Add2~2_combout  & (((\btbframes.frameblocks[2].tag [20]) # (\Add2~0_combout )))) # (!\Add2~2_combout  & (\btbframes.frameblocks[0].tag [20] & ((!\Add2~0_combout ))))

	.dataa(\btbframes.frameblocks[0].tag [20]),
	.datab(\btbframes.frameblocks[2].tag [20]),
	.datac(\Add2~2_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hF0CA;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N10
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (\Add2~0_combout  & ((\Mux8~0_combout  & (\btbframes.frameblocks[3].tag [20])) # (!\Mux8~0_combout  & ((\btbframes.frameblocks[1].tag [20]))))) # (!\Add2~0_combout  & (((\Mux8~0_combout ))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[3].tag [20]),
	.datac(\btbframes.frameblocks[1].tag [20]),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hDDA0;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N24
cycloneive_lcell_comb \does_exist~2 (
// Equation(s):
// \does_exist~2_combout  = (\Add2~42_combout  & (\Mux9~1_combout  & (\Add2~44_combout  $ (!\Mux8~1_combout )))) # (!\Add2~42_combout  & (!\Mux9~1_combout  & (\Add2~44_combout  $ (!\Mux8~1_combout ))))

	.dataa(\Add2~42_combout ),
	.datab(\Mux9~1_combout ),
	.datac(\Add2~44_combout ),
	.datad(\Mux8~1_combout ),
	.cin(gnd),
	.combout(\does_exist~2_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~2 .lut_mask = 16'h9009;
defparam \does_exist~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N16
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (\Add2~2_combout  & (((\Add2~0_combout )))) # (!\Add2~2_combout  & ((\Add2~0_combout  & (\btbframes.frameblocks[1].tag [21])) # (!\Add2~0_combout  & ((\btbframes.frameblocks[0].tag [21])))))

	.dataa(\btbframes.frameblocks[1].tag [21]),
	.datab(\btbframes.frameblocks[0].tag [21]),
	.datac(\Add2~2_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hFA0C;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N14
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (\Add2~2_combout  & ((\Mux7~0_combout  & (\btbframes.frameblocks[3].tag [21])) # (!\Mux7~0_combout  & ((\btbframes.frameblocks[2].tag [21]))))) # (!\Add2~2_combout  & (((\Mux7~0_combout ))))

	.dataa(\btbframes.frameblocks[3].tag [21]),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[2].tag [21]),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hBBC0;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N14
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (\Add2~0_combout  & (((\Add2~2_combout )))) # (!\Add2~0_combout  & ((\Add2~2_combout  & (\btbframes.frameblocks[2].tag [22])) # (!\Add2~2_combout  & ((\btbframes.frameblocks[0].tag [22])))))

	.dataa(\btbframes.frameblocks[2].tag [22]),
	.datab(\btbframes.frameblocks[0].tag [22]),
	.datac(\Add2~0_combout ),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hFA0C;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N26
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (\Mux6~0_combout  & (((\btbframes.frameblocks[3].tag [22])) # (!\Add2~0_combout ))) # (!\Mux6~0_combout  & (\Add2~0_combout  & ((\btbframes.frameblocks[1].tag [22]))))

	.dataa(\Mux6~0_combout ),
	.datab(\Add2~0_combout ),
	.datac(\btbframes.frameblocks[3].tag [22]),
	.datad(\btbframes.frameblocks[1].tag [22]),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hE6A2;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N4
cycloneive_lcell_comb \does_exist~3 (
// Equation(s):
// \does_exist~3_combout  = (\Add2~48_combout  & (\Mux6~1_combout  & (\Mux7~1_combout  $ (!\Add2~46_combout )))) # (!\Add2~48_combout  & (!\Mux6~1_combout  & (\Mux7~1_combout  $ (!\Add2~46_combout ))))

	.dataa(\Add2~48_combout ),
	.datab(\Mux7~1_combout ),
	.datac(\Add2~46_combout ),
	.datad(\Mux6~1_combout ),
	.cin(gnd),
	.combout(\does_exist~3_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~3 .lut_mask = 16'h8241;
defparam \does_exist~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N26
cycloneive_lcell_comb \does_exist~4 (
// Equation(s):
// \does_exist~4_combout  = (\does_exist~0_combout  & (\does_exist~1_combout  & (\does_exist~3_combout  & \does_exist~2_combout )))

	.dataa(\does_exist~0_combout ),
	.datab(\does_exist~1_combout ),
	.datac(\does_exist~3_combout ),
	.datad(\does_exist~2_combout ),
	.cin(gnd),
	.combout(\does_exist~4_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~4 .lut_mask = 16'h8000;
defparam \does_exist~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N8
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (\Add2~0_combout  & (((\btbframes.frameblocks[1].tag [9]) # (\Add2~2_combout )))) # (!\Add2~0_combout  & (\btbframes.frameblocks[0].tag [9] & ((!\Add2~2_combout ))))

	.dataa(\btbframes.frameblocks[0].tag [9]),
	.datab(\btbframes.frameblocks[1].tag [9]),
	.datac(\Add2~0_combout ),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hF0CA;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N26
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (\Mux19~0_combout  & (((\btbframes.frameblocks[3].tag [9]) # (!\Add2~2_combout )))) # (!\Mux19~0_combout  & (\btbframes.frameblocks[2].tag [9] & ((\Add2~2_combout ))))

	.dataa(\btbframes.frameblocks[2].tag [9]),
	.datab(\btbframes.frameblocks[3].tag [9]),
	.datac(\Mux19~0_combout ),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hCAF0;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N12
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (\Add2~2_combout  & ((\btbframes.frameblocks[2].tag [10]) # ((\Add2~0_combout )))) # (!\Add2~2_combout  & (((\btbframes.frameblocks[0].tag [10] & !\Add2~0_combout ))))

	.dataa(\Add2~2_combout ),
	.datab(\btbframes.frameblocks[2].tag [10]),
	.datac(\btbframes.frameblocks[0].tag [10]),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hAAD8;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N20
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (\Add2~0_combout  & ((\Mux18~0_combout  & ((\btbframes.frameblocks[3].tag [10]))) # (!\Mux18~0_combout  & (\btbframes.frameblocks[1].tag [10])))) # (!\Add2~0_combout  & (((\Mux18~0_combout ))))

	.dataa(\btbframes.frameblocks[1].tag [10]),
	.datab(\btbframes.frameblocks[3].tag [10]),
	.datac(\Add2~0_combout ),
	.datad(\Mux18~0_combout ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hCFA0;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N2
cycloneive_lcell_comb \does_exist~5 (
// Equation(s):
// \does_exist~5_combout  = (\Mux19~1_combout  & (\Add2~22_combout  & (\Add2~24_combout  $ (!\Mux18~1_combout )))) # (!\Mux19~1_combout  & (!\Add2~22_combout  & (\Add2~24_combout  $ (!\Mux18~1_combout ))))

	.dataa(\Mux19~1_combout ),
	.datab(\Add2~22_combout ),
	.datac(\Add2~24_combout ),
	.datad(\Mux18~1_combout ),
	.cin(gnd),
	.combout(\does_exist~5_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~5 .lut_mask = 16'h9009;
defparam \does_exist~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N14
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (\Add2~0_combout  & ((\btbframes.frameblocks[1].tag [3]) # ((\Add2~2_combout )))) # (!\Add2~0_combout  & (((\btbframes.frameblocks[0].tag [3] & !\Add2~2_combout ))))

	.dataa(\btbframes.frameblocks[1].tag [3]),
	.datab(\Add2~0_combout ),
	.datac(\btbframes.frameblocks[0].tag [3]),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hCCB8;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N26
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\Add2~2_combout  & ((\Mux25~0_combout  & ((\btbframes.frameblocks[3].tag [3]))) # (!\Mux25~0_combout  & (\btbframes.frameblocks[2].tag [3])))) # (!\Add2~2_combout  & (((\Mux25~0_combout ))))

	.dataa(\Add2~2_combout ),
	.datab(\btbframes.frameblocks[2].tag [3]),
	.datac(\btbframes.frameblocks[3].tag [3]),
	.datad(\Mux25~0_combout ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hF588;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N4
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (\Add2~0_combout  & (((\Add2~2_combout )))) # (!\Add2~0_combout  & ((\Add2~2_combout  & (\btbframes.frameblocks[2].tag [4])) # (!\Add2~2_combout  & ((\btbframes.frameblocks[0].tag [4])))))

	.dataa(\btbframes.frameblocks[2].tag [4]),
	.datab(\Add2~0_combout ),
	.datac(\btbframes.frameblocks[0].tag [4]),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hEE30;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N8
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (\Add2~0_combout  & ((\Mux24~0_combout  & ((\btbframes.frameblocks[3].tag [4]))) # (!\Mux24~0_combout  & (\btbframes.frameblocks[1].tag [4])))) # (!\Add2~0_combout  & (\Mux24~0_combout ))

	.dataa(\Add2~0_combout ),
	.datab(\Mux24~0_combout ),
	.datac(\btbframes.frameblocks[1].tag [4]),
	.datad(\btbframes.frameblocks[3].tag [4]),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hEC64;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N18
cycloneive_lcell_comb \does_exist~6 (
// Equation(s):
// \does_exist~6_combout  = (\Mux25~1_combout  & (\Add2~10_combout  & (\Mux24~1_combout  $ (!\Add2~12_combout )))) # (!\Mux25~1_combout  & (!\Add2~10_combout  & (\Mux24~1_combout  $ (!\Add2~12_combout ))))

	.dataa(\Mux25~1_combout ),
	.datab(\Add2~10_combout ),
	.datac(\Mux24~1_combout ),
	.datad(\Add2~12_combout ),
	.cin(gnd),
	.combout(\does_exist~6_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~6 .lut_mask = 16'h9009;
defparam \does_exist~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N0
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (\Add2~0_combout  & ((\btbframes.frameblocks[1].tag [5]) # ((\Add2~2_combout )))) # (!\Add2~0_combout  & (((\btbframes.frameblocks[0].tag [5] & !\Add2~2_combout ))))

	.dataa(\btbframes.frameblocks[1].tag [5]),
	.datab(\Add2~0_combout ),
	.datac(\btbframes.frameblocks[0].tag [5]),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hCCB8;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N2
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (\Add2~2_combout  & ((\Mux23~0_combout  & ((\btbframes.frameblocks[3].tag [5]))) # (!\Mux23~0_combout  & (\btbframes.frameblocks[2].tag [5])))) # (!\Add2~2_combout  & (((\Mux23~0_combout ))))

	.dataa(\btbframes.frameblocks[2].tag [5]),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[3].tag [5]),
	.datad(\Mux23~0_combout ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hF388;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N30
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (\Add2~0_combout  & (((\Add2~2_combout )))) # (!\Add2~0_combout  & ((\Add2~2_combout  & (\btbframes.frameblocks[2].tag [6])) # (!\Add2~2_combout  & ((\btbframes.frameblocks[0].tag [6])))))

	.dataa(\btbframes.frameblocks[2].tag [6]),
	.datab(\Add2~0_combout ),
	.datac(\btbframes.frameblocks[0].tag [6]),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hEE30;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N0
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (\Add2~0_combout  & ((\Mux22~0_combout  & ((\btbframes.frameblocks[3].tag [6]))) # (!\Mux22~0_combout  & (\btbframes.frameblocks[1].tag [6])))) # (!\Add2~0_combout  & (((\Mux22~0_combout ))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[1].tag [6]),
	.datac(\btbframes.frameblocks[3].tag [6]),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hF588;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N20
cycloneive_lcell_comb \does_exist~7 (
// Equation(s):
// \does_exist~7_combout  = (\Add2~14_combout  & (\Mux23~1_combout  & (\Add2~16_combout  $ (!\Mux22~1_combout )))) # (!\Add2~14_combout  & (!\Mux23~1_combout  & (\Add2~16_combout  $ (!\Mux22~1_combout ))))

	.dataa(\Add2~14_combout ),
	.datab(\Mux23~1_combout ),
	.datac(\Add2~16_combout ),
	.datad(\Mux22~1_combout ),
	.cin(gnd),
	.combout(\does_exist~7_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~7 .lut_mask = 16'h9009;
defparam \does_exist~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N6
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (\Add2~0_combout  & (((\btbframes.frameblocks[1].tag [11]) # (\Add2~2_combout )))) # (!\Add2~0_combout  & (\btbframes.frameblocks[0].tag [11] & ((!\Add2~2_combout ))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[0].tag [11]),
	.datac(\btbframes.frameblocks[1].tag [11]),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hAAE4;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N10
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (\Add2~2_combout  & ((\Mux17~0_combout  & ((\btbframes.frameblocks[3].tag [11]))) # (!\Mux17~0_combout  & (\btbframes.frameblocks[2].tag [11])))) # (!\Add2~2_combout  & (((\Mux17~0_combout ))))

	.dataa(\btbframes.frameblocks[2].tag [11]),
	.datab(\btbframes.frameblocks[3].tag [11]),
	.datac(\Add2~2_combout ),
	.datad(\Mux17~0_combout ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hCFA0;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N12
cycloneive_lcell_comb \does_exist~8 (
// Equation(s):
// \does_exist~8_combout  = (\does_exist~7_combout  & (\does_exist~6_combout  & (\Mux17~1_combout  $ (!\Add2~26_combout ))))

	.dataa(\Mux17~1_combout ),
	.datab(\does_exist~7_combout ),
	.datac(\Add2~26_combout ),
	.datad(\does_exist~6_combout ),
	.cin(gnd),
	.combout(\does_exist~8_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~8 .lut_mask = 16'h8400;
defparam \does_exist~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N18
cycloneive_lcell_comb \always3~2 (
// Equation(s):
// \always3~2_combout  = (\beq_M~q ) # (\bne_M~q )

	.dataa(gnd),
	.datab(\beq_M~q ),
	.datac(\bne_M~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\always3~2_combout ),
	.cout());
// synopsys translate_off
defparam \always3~2 .lut_mask = 16'hFCFC;
defparam \always3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N28
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (\Add2~2_combout  & (((\Add2~0_combout )))) # (!\Add2~2_combout  & ((\Add2~0_combout  & (\btbframes.frameblocks[1].tag [1])) # (!\Add2~0_combout  & ((\btbframes.frameblocks[0].tag [1])))))

	.dataa(\btbframes.frameblocks[1].tag [1]),
	.datab(\btbframes.frameblocks[0].tag [1]),
	.datac(\Add2~2_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hFA0C;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N18
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (\Add2~2_combout  & ((\Mux27~0_combout  & ((\btbframes.frameblocks[3].tag [1]))) # (!\Mux27~0_combout  & (\btbframes.frameblocks[2].tag [1])))) # (!\Add2~2_combout  & (((\Mux27~0_combout ))))

	.dataa(\btbframes.frameblocks[2].tag [1]),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[3].tag [1]),
	.datad(\Mux27~0_combout ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hF388;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N18
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (\Add2~2_combout  & ((\btbframes.frameblocks[2].tag [2]) # ((\Add2~0_combout )))) # (!\Add2~2_combout  & (((!\Add2~0_combout  & \btbframes.frameblocks[0].tag [2]))))

	.dataa(\btbframes.frameblocks[2].tag [2]),
	.datab(\Add2~2_combout ),
	.datac(\Add2~0_combout ),
	.datad(\btbframes.frameblocks[0].tag [2]),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hCBC8;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N28
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (\Add2~0_combout  & ((\Mux26~0_combout  & ((\btbframes.frameblocks[3].tag [2]))) # (!\Mux26~0_combout  & (\btbframes.frameblocks[1].tag [2])))) # (!\Add2~0_combout  & (((\Mux26~0_combout ))))

	.dataa(\btbframes.frameblocks[1].tag [2]),
	.datab(\btbframes.frameblocks[3].tag [2]),
	.datac(\Add2~0_combout ),
	.datad(\Mux26~0_combout ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hCFA0;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N28
cycloneive_lcell_comb \does_exist~9 (
// Equation(s):
// \does_exist~9_combout  = (\Add2~6_combout  & (\Mux27~1_combout  & (\Add2~8_combout  $ (!\Mux26~1_combout )))) # (!\Add2~6_combout  & (!\Mux27~1_combout  & (\Add2~8_combout  $ (!\Mux26~1_combout ))))

	.dataa(\Add2~6_combout ),
	.datab(\Mux27~1_combout ),
	.datac(\Add2~8_combout ),
	.datad(\Mux26~1_combout ),
	.cin(gnd),
	.combout(\does_exist~9_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~9 .lut_mask = 16'h9009;
defparam \does_exist~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N18
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (\Add2~0_combout  & (((\Add2~2_combout )))) # (!\Add2~0_combout  & ((\Add2~2_combout  & (\btbframes.frameblocks[2].tag [0])) # (!\Add2~2_combout  & ((\btbframes.frameblocks[0].tag [0])))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[2].tag [0]),
	.datac(\btbframes.frameblocks[0].tag [0]),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hEE50;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N30
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (\Add2~0_combout  & ((\Mux28~0_combout  & (\btbframes.frameblocks[3].tag [0])) # (!\Mux28~0_combout  & ((\btbframes.frameblocks[1].tag [0]))))) # (!\Add2~0_combout  & (((\Mux28~0_combout ))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[3].tag [0]),
	.datac(\btbframes.frameblocks[1].tag [0]),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hDDA0;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N24
cycloneive_lcell_comb \does_exist~10 (
// Equation(s):
// \does_exist~10_combout  = (\always3~2_combout  & (\does_exist~9_combout  & (\Mux28~1_combout  $ (!\Add2~4_combout ))))

	.dataa(\Mux28~1_combout ),
	.datab(\Add2~4_combout ),
	.datac(\always3~2_combout ),
	.datad(\does_exist~9_combout ),
	.cin(gnd),
	.combout(\does_exist~10_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~10 .lut_mask = 16'h9000;
defparam \does_exist~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N6
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (\Add2~2_combout  & (((\Add2~0_combout )))) # (!\Add2~2_combout  & ((\Add2~0_combout  & (\btbframes.frameblocks[1].tag [7])) # (!\Add2~0_combout  & ((\btbframes.frameblocks[0].tag [7])))))

	.dataa(\btbframes.frameblocks[1].tag [7]),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[0].tag [7]),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hEE30;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N8
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (\Add2~2_combout  & ((\Mux21~0_combout  & ((\btbframes.frameblocks[3].tag [7]))) # (!\Mux21~0_combout  & (\btbframes.frameblocks[2].tag [7])))) # (!\Add2~2_combout  & (((\Mux21~0_combout ))))

	.dataa(\Add2~2_combout ),
	.datab(\btbframes.frameblocks[2].tag [7]),
	.datac(\Mux21~0_combout ),
	.datad(\btbframes.frameblocks[3].tag [7]),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hF858;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N10
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (\Add2~0_combout  & (((\Add2~2_combout )))) # (!\Add2~0_combout  & ((\Add2~2_combout  & (\btbframes.frameblocks[2].tag [8])) # (!\Add2~2_combout  & ((\btbframes.frameblocks[0].tag [8])))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[2].tag [8]),
	.datac(\btbframes.frameblocks[0].tag [8]),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hEE50;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N10
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (\Add2~0_combout  & ((\Mux20~0_combout  & ((\btbframes.frameblocks[3].tag [8]))) # (!\Mux20~0_combout  & (\btbframes.frameblocks[1].tag [8])))) # (!\Add2~0_combout  & (((\Mux20~0_combout ))))

	.dataa(\btbframes.frameblocks[1].tag [8]),
	.datab(\btbframes.frameblocks[3].tag [8]),
	.datac(\Add2~0_combout ),
	.datad(\Mux20~0_combout ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hCFA0;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N0
cycloneive_lcell_comb \does_exist~11 (
// Equation(s):
// \does_exist~11_combout  = (\Add2~20_combout  & (\Mux20~1_combout  & (\Mux21~1_combout  $ (!\Add2~18_combout )))) # (!\Add2~20_combout  & (!\Mux20~1_combout  & (\Mux21~1_combout  $ (!\Add2~18_combout ))))

	.dataa(\Add2~20_combout ),
	.datab(\Mux21~1_combout ),
	.datac(\Add2~18_combout ),
	.datad(\Mux20~1_combout ),
	.cin(gnd),
	.combout(\does_exist~11_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~11 .lut_mask = 16'h8241;
defparam \does_exist~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N4
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (\Add2~2_combout  & ((\btbframes.frameblocks[2].tag [12]) # ((\Add2~0_combout )))) # (!\Add2~2_combout  & (((\btbframes.frameblocks[0].tag [12] & !\Add2~0_combout ))))

	.dataa(\btbframes.frameblocks[2].tag [12]),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[0].tag [12]),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hCCB8;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N24
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (\Add2~0_combout  & ((\Mux16~0_combout  & ((\btbframes.frameblocks[3].tag [12]))) # (!\Mux16~0_combout  & (\btbframes.frameblocks[1].tag [12])))) # (!\Add2~0_combout  & (((\Mux16~0_combout ))))

	.dataa(\btbframes.frameblocks[1].tag [12]),
	.datab(\Add2~0_combout ),
	.datac(\btbframes.frameblocks[3].tag [12]),
	.datad(\Mux16~0_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hF388;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N26
cycloneive_lcell_comb \does_exist~12 (
// Equation(s):
// \does_exist~12_combout  = (\does_exist~11_combout  & (\does_exist~10_combout  & (\Mux16~1_combout  $ (!\Add2~28_combout ))))

	.dataa(\Mux16~1_combout ),
	.datab(\Add2~28_combout ),
	.datac(\does_exist~11_combout ),
	.datad(\does_exist~10_combout ),
	.cin(gnd),
	.combout(\does_exist~12_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~12 .lut_mask = 16'h9000;
defparam \does_exist~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N30
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (\Add2~0_combout  & (((\btbframes.frameblocks[1].tag [13]) # (\Add2~2_combout )))) # (!\Add2~0_combout  & (\btbframes.frameblocks[0].tag [13] & ((!\Add2~2_combout ))))

	.dataa(\btbframes.frameblocks[0].tag [13]),
	.datab(\Add2~0_combout ),
	.datac(\btbframes.frameblocks[1].tag [13]),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hCCE2;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N4
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (\Add2~2_combout  & ((\Mux15~0_combout  & ((\btbframes.frameblocks[3].tag [13]))) # (!\Mux15~0_combout  & (\btbframes.frameblocks[2].tag [13])))) # (!\Add2~2_combout  & (((\Mux15~0_combout ))))

	.dataa(\Add2~2_combout ),
	.datab(\btbframes.frameblocks[2].tag [13]),
	.datac(\Mux15~0_combout ),
	.datad(\btbframes.frameblocks[3].tag [13]),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hF858;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N24
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (\Add2~2_combout  & ((\btbframes.frameblocks[2].tag [14]) # ((\Add2~0_combout )))) # (!\Add2~2_combout  & (((\btbframes.frameblocks[0].tag [14] & !\Add2~0_combout ))))

	.dataa(\btbframes.frameblocks[2].tag [14]),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[0].tag [14]),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hCCB8;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N22
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (\Add2~0_combout  & ((\Mux14~0_combout  & ((\btbframes.frameblocks[3].tag [14]))) # (!\Mux14~0_combout  & (\btbframes.frameblocks[1].tag [14])))) # (!\Add2~0_combout  & (((\Mux14~0_combout ))))

	.dataa(\btbframes.frameblocks[1].tag [14]),
	.datab(\Add2~0_combout ),
	.datac(\btbframes.frameblocks[3].tag [14]),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hF388;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N18
cycloneive_lcell_comb \does_exist~13 (
// Equation(s):
// \does_exist~13_combout  = (\Add2~30_combout  & (\Mux15~1_combout  & (\Add2~32_combout  $ (!\Mux14~1_combout )))) # (!\Add2~30_combout  & (!\Mux15~1_combout  & (\Add2~32_combout  $ (!\Mux14~1_combout ))))

	.dataa(\Add2~30_combout ),
	.datab(\Mux15~1_combout ),
	.datac(\Add2~32_combout ),
	.datad(\Mux14~1_combout ),
	.cin(gnd),
	.combout(\does_exist~13_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~13 .lut_mask = 16'h9009;
defparam \does_exist~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N20
cycloneive_lcell_comb \does_exist~14 (
// Equation(s):
// \does_exist~14_combout  = (\does_exist~13_combout  & (\does_exist~5_combout  & (\does_exist~12_combout  & \does_exist~8_combout )))

	.dataa(\does_exist~13_combout ),
	.datab(\does_exist~5_combout ),
	.datac(\does_exist~12_combout ),
	.datad(\does_exist~8_combout ),
	.cin(gnd),
	.combout(\does_exist~14_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~14 .lut_mask = 16'h8000;
defparam \does_exist~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N26
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (\Add2~2_combout  & (((\Add2~0_combout )))) # (!\Add2~2_combout  & ((\Add2~0_combout  & (\btbframes.frameblocks[1].valid~q )) # (!\Add2~0_combout  & ((\btbframes.frameblocks[0].valid~q )))))

	.dataa(\btbframes.frameblocks[1].valid~q ),
	.datab(\Add2~2_combout ),
	.datac(\Add2~0_combout ),
	.datad(\btbframes.frameblocks[0].valid~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hE3E0;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N20
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (\Mux0~0_combout  & ((\btbframes.frameblocks[3].valid~q ) # ((!\Add2~2_combout )))) # (!\Mux0~0_combout  & (((\Add2~2_combout  & \btbframes.frameblocks[2].valid~q ))))

	.dataa(\Mux0~0_combout ),
	.datab(\btbframes.frameblocks[3].valid~q ),
	.datac(\Add2~2_combout ),
	.datad(\btbframes.frameblocks[2].valid~q ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hDA8A;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N10
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (\Add2~2_combout  & (((\Add2~0_combout )))) # (!\Add2~2_combout  & ((\Add2~0_combout  & (\btbframes.frameblocks[1].tag [23])) # (!\Add2~0_combout  & ((\btbframes.frameblocks[0].tag [23])))))

	.dataa(\Add2~2_combout ),
	.datab(\btbframes.frameblocks[1].tag [23]),
	.datac(\btbframes.frameblocks[0].tag [23]),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hEE50;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N22
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (\Add2~2_combout  & ((\Mux5~0_combout  & (\btbframes.frameblocks[3].tag [23])) # (!\Mux5~0_combout  & ((\btbframes.frameblocks[2].tag [23]))))) # (!\Add2~2_combout  & (((\Mux5~0_combout ))))

	.dataa(\btbframes.frameblocks[3].tag [23]),
	.datab(\Add2~2_combout ),
	.datac(\Mux5~0_combout ),
	.datad(\btbframes.frameblocks[2].tag [23]),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hBCB0;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N10
cycloneive_lcell_comb \does_exist~15 (
// Equation(s):
// \does_exist~15_combout  = (\Mux0~1_combout  & (\does_exist~14_combout  & (\Mux5~1_combout  $ (!\Add2~50_combout ))))

	.dataa(\Mux0~1_combout ),
	.datab(\Mux5~1_combout ),
	.datac(\Add2~50_combout ),
	.datad(\does_exist~14_combout ),
	.cin(gnd),
	.combout(\does_exist~15_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~15 .lut_mask = 16'h8200;
defparam \does_exist~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N30
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (\Add2~0_combout  & (((\btbframes.frameblocks[1].tag [25]) # (\Add2~2_combout )))) # (!\Add2~0_combout  & (\btbframes.frameblocks[0].tag [25] & ((!\Add2~2_combout ))))

	.dataa(\btbframes.frameblocks[0].tag [25]),
	.datab(\btbframes.frameblocks[1].tag [25]),
	.datac(\Add2~0_combout ),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hF0CA;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N4
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (\Add2~2_combout  & ((\Mux3~0_combout  & ((\btbframes.frameblocks[3].tag [25]))) # (!\Mux3~0_combout  & (\btbframes.frameblocks[2].tag [25])))) # (!\Add2~2_combout  & (((\Mux3~0_combout ))))

	.dataa(\Add2~2_combout ),
	.datab(\btbframes.frameblocks[2].tag [25]),
	.datac(\Mux3~0_combout ),
	.datad(\btbframes.frameblocks[3].tag [25]),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hF858;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N6
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (\Add2~2_combout  & (((\btbframes.frameblocks[2].tag [24]) # (\Add2~0_combout )))) # (!\Add2~2_combout  & (\btbframes.frameblocks[0].tag [24] & ((!\Add2~0_combout ))))

	.dataa(\btbframes.frameblocks[0].tag [24]),
	.datab(\btbframes.frameblocks[2].tag [24]),
	.datac(\Add2~2_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hF0CA;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N6
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (\Mux4~0_combout  & ((\btbframes.frameblocks[3].tag [24]) # ((!\Add2~0_combout )))) # (!\Mux4~0_combout  & (((\Add2~0_combout  & \btbframes.frameblocks[1].tag [24]))))

	.dataa(\Mux4~0_combout ),
	.datab(\btbframes.frameblocks[3].tag [24]),
	.datac(\Add2~0_combout ),
	.datad(\btbframes.frameblocks[1].tag [24]),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hDA8A;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N18
cycloneive_lcell_comb \does_exist~16 (
// Equation(s):
// \does_exist~16_combout  = (\Add2~54_combout  & (\Mux3~1_combout  & (\Add2~52_combout  $ (!\Mux4~1_combout )))) # (!\Add2~54_combout  & (!\Mux3~1_combout  & (\Add2~52_combout  $ (!\Mux4~1_combout ))))

	.dataa(\Add2~54_combout ),
	.datab(\Mux3~1_combout ),
	.datac(\Add2~52_combout ),
	.datad(\Mux4~1_combout ),
	.cin(gnd),
	.combout(\does_exist~16_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~16 .lut_mask = 16'h9009;
defparam \does_exist~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N22
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (\Add2~0_combout  & ((\btbframes.frameblocks[1].tag [27]) # ((\Add2~2_combout )))) # (!\Add2~0_combout  & (((\btbframes.frameblocks[0].tag [27] & !\Add2~2_combout ))))

	.dataa(\Add2~0_combout ),
	.datab(\btbframes.frameblocks[1].tag [27]),
	.datac(\btbframes.frameblocks[0].tag [27]),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hAAD8;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N0
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (\Mux1~0_combout  & (((\btbframes.frameblocks[3].tag [27]) # (!\Add2~2_combout )))) # (!\Mux1~0_combout  & (\btbframes.frameblocks[2].tag [27] & ((\Add2~2_combout ))))

	.dataa(\btbframes.frameblocks[2].tag [27]),
	.datab(\btbframes.frameblocks[3].tag [27]),
	.datac(\Mux1~0_combout ),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hCAF0;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N12
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (\Add2~0_combout  & (\Add2~2_combout )) # (!\Add2~0_combout  & ((\Add2~2_combout  & ((\btbframes.frameblocks[2].tag [26]))) # (!\Add2~2_combout  & (\btbframes.frameblocks[0].tag [26]))))

	.dataa(\Add2~0_combout ),
	.datab(\Add2~2_combout ),
	.datac(\btbframes.frameblocks[0].tag [26]),
	.datad(\btbframes.frameblocks[2].tag [26]),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hDC98;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N24
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (\Add2~0_combout  & ((\Mux2~0_combout  & (\btbframes.frameblocks[3].tag [26])) # (!\Mux2~0_combout  & ((\btbframes.frameblocks[1].tag [26]))))) # (!\Add2~0_combout  & (((\Mux2~0_combout ))))

	.dataa(\btbframes.frameblocks[3].tag [26]),
	.datab(\Add2~0_combout ),
	.datac(\btbframes.frameblocks[1].tag [26]),
	.datad(\Mux2~0_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hBBC0;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N2
cycloneive_lcell_comb \does_exist~17 (
// Equation(s):
// \does_exist~17_combout  = (\Add2~58_combout  & (\Mux1~1_combout  & (\Mux2~1_combout  $ (!\Add2~56_combout )))) # (!\Add2~58_combout  & (!\Mux1~1_combout  & (\Mux2~1_combout  $ (!\Add2~56_combout ))))

	.dataa(\Add2~58_combout ),
	.datab(\Mux1~1_combout ),
	.datac(\Mux2~1_combout ),
	.datad(\Add2~56_combout ),
	.cin(gnd),
	.combout(\does_exist~17_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~17 .lut_mask = 16'h9009;
defparam \does_exist~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N0
cycloneive_lcell_comb \does_exist~18 (
// Equation(s):
// \does_exist~18_combout  = (\does_exist~4_combout  & (\does_exist~16_combout  & (\does_exist~17_combout  & \does_exist~15_combout )))

	.dataa(\does_exist~4_combout ),
	.datab(\does_exist~16_combout ),
	.datac(\does_exist~17_combout ),
	.datad(\does_exist~15_combout ),
	.cin(gnd),
	.combout(\does_exist~18_combout ),
	.cout());
// synopsys translate_off
defparam \does_exist~18 .lut_mask = 16'h8000;
defparam \does_exist~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N6
cycloneive_lcell_comb \btbframes.frameblocks[2].tag[27]~2 (
// Equation(s):
// \btbframes.frameblocks[2].tag[27]~2_combout  = (\btbframes.frameblocks[2].tag[27]~3_combout  & (\Decoder0~0_combout  & (iwait & !\does_exist~18_combout )))

	.dataa(\btbframes.frameblocks[2].tag[27]~3_combout ),
	.datab(\Decoder0~0_combout ),
	.datac(iwait),
	.datad(\does_exist~18_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].tag[27]~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[27]~2 .lut_mask = 16'h0080;
defparam \btbframes.frameblocks[2].tag[27]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N22
cycloneive_lcell_comb \Decoder0~1 (
// Equation(s):
// \Decoder0~1_combout  = (!\Add2~2_combout  & \Add2~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~2_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~1 .lut_mask = 16'h0F00;
defparam \Decoder0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N4
cycloneive_lcell_comb \btbframes.frameblocks[1].tag[27]~2 (
// Equation(s):
// \btbframes.frameblocks[1].tag[27]~2_combout  = (\btbframes.frameblocks[2].tag[27]~3_combout  & (\Decoder0~1_combout  & (iwait & !\does_exist~18_combout )))

	.dataa(\btbframes.frameblocks[2].tag[27]~3_combout ),
	.datab(\Decoder0~1_combout ),
	.datac(iwait),
	.datad(\does_exist~18_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].tag[27]~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[27]~2 .lut_mask = 16'h0080;
defparam \btbframes.frameblocks[1].tag[27]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N18
cycloneive_lcell_comb \btbframes.frameblocks[0].tag[27]~2 (
// Equation(s):
// \btbframes.frameblocks[0].tag[27]~2_combout  = (\btbframes.frameblocks[0].tag[27]~3_combout  & (!\Add2~0_combout  & (iwait & !\does_exist~18_combout )))

	.dataa(\btbframes.frameblocks[0].tag[27]~3_combout ),
	.datab(\Add2~0_combout ),
	.datac(iwait),
	.datad(\does_exist~18_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].tag[27]~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[27]~2 .lut_mask = 16'h0020;
defparam \btbframes.frameblocks[0].tag[27]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N8
cycloneive_lcell_comb \Decoder0~2 (
// Equation(s):
// \Decoder0~2_combout  = (\Add2~0_combout  & \Add2~2_combout )

	.dataa(gnd),
	.datab(\Add2~0_combout ),
	.datac(gnd),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~2 .lut_mask = 16'hCC00;
defparam \Decoder0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N30
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[27]~2 (
// Equation(s):
// \btbframes.frameblocks[3].tag[27]~2_combout  = (\btbframes.frameblocks[2].tag[27]~3_combout  & (\Decoder0~2_combout  & (iwait & !\does_exist~18_combout )))

	.dataa(\btbframes.frameblocks[2].tag[27]~3_combout ),
	.datab(\Decoder0~2_combout ),
	.datac(iwait),
	.datad(\does_exist~18_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[27]~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[27]~2 .lut_mask = 16'h0080;
defparam \btbframes.frameblocks[3].tag[27]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N18
cycloneive_lcell_comb \rdata1_M~32 (
// Equation(s):
// \rdata1_M~32_combout  = (fuifforward_A_0 & (\regWrite_M~q  & (!Equal31 & \jr_EX~q )))

	.dataa(\FORWARDING_UNIT|fuif.forward_A[0]~2_combout ),
	.datab(\regWrite_M~q ),
	.datac(\FORWARDING_UNIT|Equal3~1_combout ),
	.datad(\jr_EX~q ),
	.cin(gnd),
	.combout(\rdata1_M~32_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M~32 .lut_mask = 16'h0800;
defparam \rdata1_M~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N28
cycloneive_lcell_comb \rdata1_M~33 (
// Equation(s):
// \rdata1_M~33_combout  = (\jr_EX~q  & (fuifforward_A_11 & !fuifforward_A_01))

	.dataa(gnd),
	.datab(\jr_EX~q ),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\rdata1_M~33_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_M~33 .lut_mask = 16'h00C0;
defparam \rdata1_M~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N13
dffeas \pc_plus_4_EX[1] (
	.clk(CLK),
	.d(\pc_plus_4_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[1]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[1] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N26
cycloneive_lcell_comb \btbframes.frameblocks[0].valid~0 (
// Equation(s):
// \btbframes.frameblocks[0].valid~0_combout  = (\btbframes.frameblocks[0].valid~q ) # ((!\Add2~2_combout  & (\always3~3_combout  & !\Add2~0_combout )))

	.dataa(\Add2~2_combout ),
	.datab(\always3~3_combout ),
	.datac(\btbframes.frameblocks[0].valid~q ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].valid~0_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].valid~0 .lut_mask = 16'hF0F4;
defparam \btbframes.frameblocks[0].valid~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N8
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (\Add2~0_combout  & (((\Add2~2_combout )))) # (!\Add2~0_combout  & ((\Add2~2_combout  & (\btbframes.frameblocks[2].curr_state [1])) # (!\Add2~2_combout  & ((\btbframes.frameblocks[0].curr_state [1])))))

	.dataa(\btbframes.frameblocks[2].curr_state [1]),
	.datab(\Add2~0_combout ),
	.datac(\btbframes.frameblocks[0].curr_state [1]),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hEE30;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N26
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (\Mux29~0_combout  & ((\btbframes.frameblocks[3].curr_state [1]) # ((!\Add2~0_combout )))) # (!\Mux29~0_combout  & (((\btbframes.frameblocks[1].curr_state [1] & \Add2~0_combout ))))

	.dataa(\btbframes.frameblocks[3].curr_state [1]),
	.datab(\btbframes.frameblocks[1].curr_state [1]),
	.datac(\Mux29~0_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hACF0;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N17
dffeas \btbframes.frameblocks[2].curr_state[0] (
	.clk(CLK),
	.d(\btbframes.frameblocks[2].curr_state[0]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[2].curr_state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[2].curr_state[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[2].curr_state[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N11
dffeas \btbframes.frameblocks[1].curr_state[0] (
	.clk(CLK),
	.d(\btbframes.frameblocks[1].curr_state[0]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[1].curr_state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[1].curr_state[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[1].curr_state[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N21
dffeas \btbframes.frameblocks[0].curr_state[0] (
	.clk(CLK),
	.d(\btbframes.frameblocks[0].curr_state[0]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[0].curr_state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[0].curr_state[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[0].curr_state[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N30
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (\Add2~2_combout  & (((\Add2~0_combout )))) # (!\Add2~2_combout  & ((\Add2~0_combout  & (!\btbframes.frameblocks[1].curr_state [0])) # (!\Add2~0_combout  & ((!\btbframes.frameblocks[0].curr_state [0])))))

	.dataa(\btbframes.frameblocks[1].curr_state [0]),
	.datab(\btbframes.frameblocks[0].curr_state [0]),
	.datac(\Add2~2_combout ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hF503;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y40_N13
dffeas \btbframes.frameblocks[3].curr_state[0] (
	.clk(CLK),
	.d(\btbframes.frameblocks[3].curr_state[0]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\btbframes.frameblocks[3].curr_state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \btbframes.frameblocks[3].curr_state[0] .is_wysiwyg = "true";
defparam \btbframes.frameblocks[3].curr_state[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N14
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (\Mux30~0_combout  & (((!\Add2~2_combout )) # (!\btbframes.frameblocks[3].curr_state [0]))) # (!\Mux30~0_combout  & (((!\btbframes.frameblocks[2].curr_state [0] & \Add2~2_combout ))))

	.dataa(\btbframes.frameblocks[3].curr_state [0]),
	.datab(\btbframes.frameblocks[2].curr_state [0]),
	.datac(\Mux30~0_combout ),
	.datad(\Add2~2_combout ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'h53F0;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N24
cycloneive_lcell_comb \btbframes~0 (
// Equation(s):
// \btbframes~0_combout  = (iwait & ((\does_exist~18_combout  & ((\branch_taken~0_combout ))) # (!\does_exist~18_combout  & (\always3~2_combout ))))

	.dataa(\always3~2_combout ),
	.datab(iwait),
	.datac(\does_exist~18_combout ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\btbframes~0_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes~0 .lut_mask = 16'hC808;
defparam \btbframes~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N18
cycloneive_lcell_comb \btbframes~1 (
// Equation(s):
// \btbframes~1_combout  = (\Mux29~1_combout  & (((!\Mux30~1_combout  & !\always3~3_combout )) # (!\btbframes~0_combout ))) # (!\Mux29~1_combout  & (!\Mux30~1_combout  & ((!\btbframes~0_combout ))))

	.dataa(\Mux29~1_combout ),
	.datab(\Mux30~1_combout ),
	.datac(\always3~3_combout ),
	.datad(\btbframes~0_combout ),
	.cin(gnd),
	.combout(\btbframes~1_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes~1 .lut_mask = 16'h02BB;
defparam \btbframes~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N12
cycloneive_lcell_comb \btbframes.frameblocks[2].curr_state[0]~0 (
// Equation(s):
// \btbframes.frameblocks[2].curr_state[0]~0_combout  = (\branch_taken~0_combout  & ((\Mux29~1_combout ) # (!\Mux30~1_combout )))

	.dataa(gnd),
	.datab(\branch_taken~0_combout ),
	.datac(\Mux29~1_combout ),
	.datad(\Mux30~1_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].curr_state[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].curr_state[0]~0 .lut_mask = 16'hC0CC;
defparam \btbframes.frameblocks[2].curr_state[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N26
cycloneive_lcell_comb \btbframes.frameblocks[2].curr_state[0]~1 (
// Equation(s):
// \btbframes.frameblocks[2].curr_state[0]~1_combout  = (iwait & ((\does_exist~18_combout  & (\btbframes.frameblocks[2].curr_state[0]~0_combout )) # (!\does_exist~18_combout  & ((\always3~2_combout )))))

	.dataa(\btbframes.frameblocks[2].curr_state[0]~0_combout ),
	.datab(\always3~2_combout ),
	.datac(iwait),
	.datad(\does_exist~18_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].curr_state[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].curr_state[0]~1 .lut_mask = 16'hA0C0;
defparam \btbframes.frameblocks[2].curr_state[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N8
cycloneive_lcell_comb \btbframes.frameblocks[1].curr_state[1]~0 (
// Equation(s):
// \btbframes.frameblocks[1].curr_state[1]~0_combout  = (\Mux30~1_combout ) # (!\Mux29~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux29~1_combout ),
	.datad(\Mux30~1_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].curr_state[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].curr_state[1]~0 .lut_mask = 16'hFF0F;
defparam \btbframes.frameblocks[1].curr_state[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N6
cycloneive_lcell_comb \btbframes.frameblocks[1].curr_state[1]~1 (
// Equation(s):
// \btbframes.frameblocks[1].curr_state[1]~1_combout  = (\btbframes.frameblocks[1].curr_state[1]~0_combout  & (!\branch_taken~0_combout  & (iwait & \does_exist~18_combout )))

	.dataa(\btbframes.frameblocks[1].curr_state[1]~0_combout ),
	.datab(\branch_taken~0_combout ),
	.datac(iwait),
	.datad(\does_exist~18_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].curr_state[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].curr_state[1]~1 .lut_mask = 16'h2000;
defparam \btbframes.frameblocks[1].curr_state[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N28
cycloneive_lcell_comb \btbframes.frameblocks[2].curr_state[1]~2 (
// Equation(s):
// \btbframes.frameblocks[2].curr_state[1]~2_combout  = (\nRST~input_o  & ((\btbframes.frameblocks[2].curr_state[0]~1_combout ) # (\btbframes.frameblocks[1].curr_state[1]~1_combout )))

	.dataa(gnd),
	.datab(nRST),
	.datac(\btbframes.frameblocks[2].curr_state[0]~1_combout ),
	.datad(\btbframes.frameblocks[1].curr_state[1]~1_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].curr_state[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].curr_state[1]~2 .lut_mask = 16'hCCC0;
defparam \btbframes.frameblocks[2].curr_state[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N4
cycloneive_lcell_comb \btbframes.frameblocks[1].curr_state[1]~2 (
// Equation(s):
// \btbframes.frameblocks[1].curr_state[1]~2_combout  = (\Decoder0~1_combout  & ((\btbframes.frameblocks[2].curr_state[1]~2_combout  & (\btbframes~1_combout )) # (!\btbframes.frameblocks[2].curr_state[1]~2_combout  & ((\btbframes.frameblocks[1].curr_state 
// [1]))))) # (!\Decoder0~1_combout  & (((\btbframes.frameblocks[1].curr_state [1]))))

	.dataa(\Decoder0~1_combout ),
	.datab(\btbframes~1_combout ),
	.datac(\btbframes.frameblocks[1].curr_state [1]),
	.datad(\btbframes.frameblocks[2].curr_state[1]~2_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].curr_state[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].curr_state[1]~2 .lut_mask = 16'hD8F0;
defparam \btbframes.frameblocks[1].curr_state[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N6
cycloneive_lcell_comb \btbframes.frameblocks[2].curr_state[1]~3 (
// Equation(s):
// \btbframes.frameblocks[2].curr_state[1]~3_combout  = (\Decoder0~0_combout  & ((\btbframes.frameblocks[2].curr_state[1]~2_combout  & (\btbframes~1_combout )) # (!\btbframes.frameblocks[2].curr_state[1]~2_combout  & ((\btbframes.frameblocks[2].curr_state 
// [1]))))) # (!\Decoder0~0_combout  & (((\btbframes.frameblocks[2].curr_state [1]))))

	.dataa(\Decoder0~0_combout ),
	.datab(\btbframes~1_combout ),
	.datac(\btbframes.frameblocks[2].curr_state [1]),
	.datad(\btbframes.frameblocks[2].curr_state[1]~2_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].curr_state[1]~3_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].curr_state[1]~3 .lut_mask = 16'hD8F0;
defparam \btbframes.frameblocks[2].curr_state[1]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N22
cycloneive_lcell_comb \btbframes.frameblocks[0].curr_state[1]~0 (
// Equation(s):
// \btbframes.frameblocks[0].curr_state[1]~0_combout  = (\nRST~input_o  & !\Add2~0_combout )

	.dataa(gnd),
	.datab(nRST),
	.datac(\Add2~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].curr_state[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].curr_state[1]~0 .lut_mask = 16'h0C0C;
defparam \btbframes.frameblocks[0].curr_state[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N4
cycloneive_lcell_comb \btbframes.frameblocks[0].curr_state[1]~1 (
// Equation(s):
// \btbframes.frameblocks[0].curr_state[1]~1_combout  = (!\Add2~2_combout  & (\btbframes.frameblocks[0].curr_state[1]~0_combout  & ((\btbframes.frameblocks[2].curr_state[0]~1_combout ) # (\btbframes.frameblocks[1].curr_state[1]~1_combout ))))

	.dataa(\Add2~2_combout ),
	.datab(\btbframes.frameblocks[0].curr_state[1]~0_combout ),
	.datac(\btbframes.frameblocks[2].curr_state[0]~1_combout ),
	.datad(\btbframes.frameblocks[1].curr_state[1]~1_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].curr_state[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].curr_state[1]~1 .lut_mask = 16'h4440;
defparam \btbframes.frameblocks[0].curr_state[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N28
cycloneive_lcell_comb \btbframes.frameblocks[0].curr_state[1]~2 (
// Equation(s):
// \btbframes.frameblocks[0].curr_state[1]~2_combout  = (\btbframes.frameblocks[0].curr_state[1]~1_combout  & (\btbframes~1_combout )) # (!\btbframes.frameblocks[0].curr_state[1]~1_combout  & ((\btbframes.frameblocks[0].curr_state [1])))

	.dataa(gnd),
	.datab(\btbframes~1_combout ),
	.datac(\btbframes.frameblocks[0].curr_state [1]),
	.datad(\btbframes.frameblocks[0].curr_state[1]~1_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].curr_state[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].curr_state[1]~2 .lut_mask = 16'hCCF0;
defparam \btbframes.frameblocks[0].curr_state[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N22
cycloneive_lcell_comb \btbframes.frameblocks[3].curr_state[1]~0 (
// Equation(s):
// \btbframes.frameblocks[3].curr_state[1]~0_combout  = (\Decoder0~2_combout  & ((\btbframes.frameblocks[2].curr_state[1]~2_combout  & (\btbframes~1_combout )) # (!\btbframes.frameblocks[2].curr_state[1]~2_combout  & ((\btbframes.frameblocks[3].curr_state 
// [1]))))) # (!\Decoder0~2_combout  & (((\btbframes.frameblocks[3].curr_state [1]))))

	.dataa(\Decoder0~2_combout ),
	.datab(\btbframes~1_combout ),
	.datac(\btbframes.frameblocks[3].curr_state [1]),
	.datad(\btbframes.frameblocks[2].curr_state[1]~2_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].curr_state[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].curr_state[1]~0 .lut_mask = 16'hD8F0;
defparam \btbframes.frameblocks[3].curr_state[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N21
dffeas \pc_plus_4_EX[8] (
	.clk(CLK),
	.d(\pc_plus_4_EX~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[8]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[8] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N15
dffeas \pc_plus_4_EX[12] (
	.clk(CLK),
	.d(\pc_plus_4_EX~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[12]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[12] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N3
dffeas \pc_plus_4_EX[15] (
	.clk(CLK),
	.d(\pc_plus_4_EX~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[15]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[15] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N7
dffeas \pc_plus_4_EX[14] (
	.clk(CLK),
	.d(\pc_plus_4_EX~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[14]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[14] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N9
dffeas \pc_plus_4_EX[16] (
	.clk(CLK),
	.d(\pc_plus_4_EX~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[16]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[16] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N6
cycloneive_lcell_comb \pc_plus_4_M~17 (
// Equation(s):
// \pc_plus_4_M~17_combout  = (pc_plus_4_EX[16] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[16]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~17_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~17 .lut_mask = 16'h00CC;
defparam \pc_plus_4_M~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N17
dffeas \pc_plus_4_EX[18] (
	.clk(CLK),
	.d(\pc_plus_4_EX~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[18]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[18] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N0
cycloneive_lcell_comb \pc_plus_4_M~19 (
// Equation(s):
// \pc_plus_4_M~19_combout  = (pc_plus_4_EX[18] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[18]),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_plus_4_M~19_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~19 .lut_mask = 16'h0C0C;
defparam \pc_plus_4_M~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N18
cycloneive_lcell_comb \instruction_M~0 (
// Equation(s):
// \instruction_M~0_combout  = (instruction_EX[17] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(instruction_EX[17]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\instruction_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_M~0 .lut_mask = 16'h00CC;
defparam \instruction_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N30
cycloneive_lcell_comb \instruction_M~1 (
// Equation(s):
// \instruction_M~1_combout  = (!\wsel_M~0_combout  & instruction_EX[16])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(instruction_EX[16]),
	.cin(gnd),
	.combout(\instruction_M~1_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_M~1 .lut_mask = 16'h0F00;
defparam \instruction_M~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N1
dffeas \pc_plus_4_EX[21] (
	.clk(CLK),
	.d(\pc_plus_4_EX~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[21]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[21] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N28
cycloneive_lcell_comb \pc_plus_4_M~20 (
// Equation(s):
// \pc_plus_4_M~20_combout  = (pc_plus_4_EX[21] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[21]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~20_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~20 .lut_mask = 16'h00CC;
defparam \pc_plus_4_M~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N26
cycloneive_lcell_comb \instruction_M~2 (
// Equation(s):
// \instruction_M~2_combout  = (!\wsel_M~0_combout  & instruction_EX[19])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(instruction_EX[19]),
	.cin(gnd),
	.combout(\instruction_M~2_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_M~2 .lut_mask = 16'h0F00;
defparam \instruction_M~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N30
cycloneive_lcell_comb \instruction_M~3 (
// Equation(s):
// \instruction_M~3_combout  = (!\wsel_M~0_combout  & instruction_EX[18])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(instruction_EX[18]),
	.cin(gnd),
	.combout(\instruction_M~3_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_M~3 .lut_mask = 16'h0F00;
defparam \instruction_M~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N23
dffeas \pc_plus_4_EX[22] (
	.clk(CLK),
	.d(\pc_plus_4_EX~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[22]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[22] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N4
cycloneive_lcell_comb \instruction_M~4 (
// Equation(s):
// \instruction_M~4_combout  = (instruction_EX[21] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(instruction_EX[21]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\instruction_M~4_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_M~4 .lut_mask = 16'h00CC;
defparam \instruction_M~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N22
cycloneive_lcell_comb \instruction_M~5 (
// Equation(s):
// \instruction_M~5_combout  = (instruction_EX[20] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(instruction_EX[20]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\instruction_M~5_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_M~5 .lut_mask = 16'h00CC;
defparam \instruction_M~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N12
cycloneive_lcell_comb \instruction_M~6 (
// Equation(s):
// \instruction_M~6_combout  = (instruction_EX[23] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(instruction_EX[23]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\instruction_M~6_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_M~6 .lut_mask = 16'h00CC;
defparam \instruction_M~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N28
cycloneive_lcell_comb \instruction_M~7 (
// Equation(s):
// \instruction_M~7_combout  = (instruction_EX[22] & !\wsel_M~0_combout )

	.dataa(instruction_EX[22]),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\instruction_M~7_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_M~7 .lut_mask = 16'h0A0A;
defparam \instruction_M~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N0
cycloneive_lcell_comb \instruction_M~8 (
// Equation(s):
// \instruction_M~8_combout  = (instruction_EX[25] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(instruction_EX[25]),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\instruction_M~8_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_M~8 .lut_mask = 16'h00F0;
defparam \instruction_M~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N22
cycloneive_lcell_comb \instruction_M~9 (
// Equation(s):
// \instruction_M~9_combout  = (instruction_EX[24] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(instruction_EX[24]),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\instruction_M~9_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_M~9 .lut_mask = 16'h0C0C;
defparam \instruction_M~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N25
dffeas \pc_plus_4_EX[29] (
	.clk(CLK),
	.d(\pc_plus_4_EX~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[29]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[29] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N31
dffeas \pc_plus_4_EX[28] (
	.clk(CLK),
	.d(\pc_plus_4_EX~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[28]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[28] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N22
cycloneive_lcell_comb \pc_plus_4_M~29 (
// Equation(s):
// \pc_plus_4_M~29_combout  = (pc_plus_4_EX[28] & !\wsel_M~0_combout )

	.dataa(pc_plus_4_EX[28]),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_plus_4_M~29_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~29 .lut_mask = 16'h0A0A;
defparam \pc_plus_4_M~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N12
cycloneive_lcell_comb \sw_forwarding_output~29 (
// Equation(s):
// \sw_forwarding_output~29_combout  = (!\lui_M~q  & porto_M_2)

	.dataa(gnd),
	.datab(gnd),
	.datac(\lui_M~q ),
	.datad(porto_M_2),
	.cin(gnd),
	.combout(\sw_forwarding_output~29_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~29 .lut_mask = 16'h0F00;
defparam \sw_forwarding_output~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N26
cycloneive_lcell_comb \sw_forwarding_output~31 (
// Equation(s):
// \sw_forwarding_output~31_combout  = (!\lui_M~q  & porto_M_4)

	.dataa(\lui_M~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(porto_M_4),
	.cin(gnd),
	.combout(\sw_forwarding_output~31_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~31 .lut_mask = 16'h5500;
defparam \sw_forwarding_output~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N12
cycloneive_lcell_comb \cu_halt_EX~0 (
// Equation(s):
// \cu_halt_EX~0_combout  = (\branch_or_jump~1_combout  & Decoder11)

	.dataa(gnd),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\CONTROL_UNIT|Decoder1~1_combout ),
	.cin(gnd),
	.combout(\cu_halt_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \cu_halt_EX~0 .lut_mask = 16'hF000;
defparam \cu_halt_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N11
dffeas predicted_D(
	.clk(CLK),
	.d(\predicted_D~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\predicted_D~q ),
	.prn(vcc));
// synopsys translate_off
defparam predicted_D.is_wysiwyg = "true";
defparam predicted_D.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N24
cycloneive_lcell_comb \predicted_EX~0 (
// Equation(s):
// \predicted_EX~0_combout  = (\predicted_D~q  & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\predicted_D~q ),
	.datab(\branch_or_jump~2_combout ),
	.datac(\branch_taken~0_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\predicted_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \predicted_EX~0 .lut_mask = 16'h8008;
defparam \predicted_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N16
cycloneive_lcell_comb \jr_EX~0 (
// Equation(s):
// \jr_EX~0_combout  = (\branch_or_jump~1_combout  & (!Decoder0 & Equal31))

	.dataa(\branch_or_jump~1_combout ),
	.datab(\CONTROL_UNIT|Decoder0~1_combout ),
	.datac(\CONTROL_UNIT|Equal3~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\jr_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \jr_EX~0 .lut_mask = 16'h2020;
defparam \jr_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N2
cycloneive_lcell_comb \op_D~0 (
// Equation(s):
// \op_D~0_combout  = (iwait & (((ramiframload_31)))) # (!iwait & (instruction_D[31] & (!\always2~2_combout )))

	.dataa(instruction_D[31]),
	.datab(\always2~2_combout ),
	.datac(\dpif.dmemload [31]),
	.datad(iwait),
	.cin(gnd),
	.combout(\op_D~0_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~0 .lut_mask = 16'hF022;
defparam \op_D~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N4
cycloneive_lcell_comb \op_D~1 (
// Equation(s):
// \op_D~1_combout  = (!\op_D~0_combout ) # (!\branch_or_jump~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\op_D~0_combout ),
	.cin(gnd),
	.combout(\op_D~1_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~1 .lut_mask = 16'h0FFF;
defparam \op_D~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N2
cycloneive_lcell_comb \op_D~2 (
// Equation(s):
// \op_D~2_combout  = (instruction_D[30] & (dhit & (fuifbubble_lw_f & always1)))

	.dataa(instruction_D[30]),
	.datab(dhit),
	.datac(\FORWARDING_UNIT|fuif.bubble_lw_f~2_combout ),
	.datad(always1),
	.cin(gnd),
	.combout(\op_D~2_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~2 .lut_mask = 16'h8000;
defparam \op_D~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N28
cycloneive_lcell_comb \op_D~3 (
// Equation(s):
// \op_D~3_combout  = ((!\op_D~2_combout  & ((!ramiframload_30) # (!iwait)))) # (!\branch_or_jump~1_combout )

	.dataa(iwait),
	.datab(\op_D~2_combout ),
	.datac(\branch_or_jump~1_combout ),
	.datad(\dpif.dmemload [30]),
	.cin(gnd),
	.combout(\op_D~3_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~3 .lut_mask = 16'h1F3F;
defparam \op_D~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N12
cycloneive_lcell_comb \op_D~4 (
// Equation(s):
// \op_D~4_combout  = (iwait & (((ramiframload_29)))) # (!iwait & (instruction_D[29] & (!\always2~2_combout )))

	.dataa(iwait),
	.datab(instruction_D[29]),
	.datac(\always2~2_combout ),
	.datad(\dpif.dmemload [29]),
	.cin(gnd),
	.combout(\op_D~4_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~4 .lut_mask = 16'hAE04;
defparam \op_D~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N14
cycloneive_lcell_comb \op_D~5 (
// Equation(s):
// \op_D~5_combout  = (!\op_D~4_combout ) # (!\branch_or_jump~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\op_D~4_combout ),
	.cin(gnd),
	.combout(\op_D~5_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~5 .lut_mask = 16'h0FFF;
defparam \op_D~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N24
cycloneive_lcell_comb \op_D~6 (
// Equation(s):
// \op_D~6_combout  = (fuifbubble_lw_f & (dhit & (instruction_D[28] & always1)))

	.dataa(\FORWARDING_UNIT|fuif.bubble_lw_f~2_combout ),
	.datab(dhit),
	.datac(instruction_D[28]),
	.datad(always1),
	.cin(gnd),
	.combout(\op_D~6_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~6 .lut_mask = 16'h8000;
defparam \op_D~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N26
cycloneive_lcell_comb \op_D~7 (
// Equation(s):
// \op_D~7_combout  = ((!\op_D~6_combout  & ((!iwait) # (!ramiframload_28)))) # (!\branch_or_jump~1_combout )

	.dataa(\op_D~6_combout ),
	.datab(\branch_or_jump~1_combout ),
	.datac(\dpif.dmemload [28]),
	.datad(iwait),
	.cin(gnd),
	.combout(\op_D~7_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~7 .lut_mask = 16'h3777;
defparam \op_D~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N10
cycloneive_lcell_comb \op_D~8 (
// Equation(s):
// \op_D~8_combout  = (iwait & (((ramiframload_27)))) # (!iwait & (instruction_D[27] & (!\always2~2_combout )))

	.dataa(iwait),
	.datab(instruction_D[27]),
	.datac(\always2~2_combout ),
	.datad(\dpif.dmemload [27]),
	.cin(gnd),
	.combout(\op_D~8_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~8 .lut_mask = 16'hAE04;
defparam \op_D~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N8
cycloneive_lcell_comb \op_D~9 (
// Equation(s):
// \op_D~9_combout  = (!\op_D~8_combout ) # (!\branch_or_jump~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\op_D~8_combout ),
	.cin(gnd),
	.combout(\op_D~9_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~9 .lut_mask = 16'h0FFF;
defparam \op_D~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N24
cycloneive_lcell_comb \op_D~10 (
// Equation(s):
// \op_D~10_combout  = (iwait & (((ramiframload_26)))) # (!iwait & (instruction_D[26] & (!\always2~2_combout )))

	.dataa(iwait),
	.datab(instruction_D[26]),
	.datac(\always2~2_combout ),
	.datad(\dpif.dmemload [26]),
	.cin(gnd),
	.combout(\op_D~10_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~10 .lut_mask = 16'hAE04;
defparam \op_D~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N6
cycloneive_lcell_comb \op_D~11 (
// Equation(s):
// \op_D~11_combout  = (!\op_D~10_combout ) # (!\branch_or_jump~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\op_D~10_combout ),
	.cin(gnd),
	.combout(\op_D~11_combout ),
	.cout());
// synopsys translate_off
defparam \op_D~11 .lut_mask = 16'h0FFF;
defparam \op_D~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N26
cycloneive_lcell_comb \RegDst_EX~0 (
// Equation(s):
// \RegDst_EX~0_combout  = (\branch_or_jump~1_combout  & Equal31)

	.dataa(gnd),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\CONTROL_UNIT|Equal3~2_combout ),
	.cin(gnd),
	.combout(\RegDst_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \RegDst_EX~0 .lut_mask = 16'hF000;
defparam \RegDst_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N28
cycloneive_lcell_comb \RegWrite_EX~0 (
// Equation(s):
// \RegWrite_EX~0_combout  = (instruction_D[29]) # ((instruction_D[26] & instruction_D[27]))

	.dataa(instruction_D[26]),
	.datab(gnd),
	.datac(instruction_D[29]),
	.datad(instruction_D[27]),
	.cin(gnd),
	.combout(\RegWrite_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \RegWrite_EX~0 .lut_mask = 16'hFAF0;
defparam \RegWrite_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N22
cycloneive_lcell_comb \RegWrite_EX~1 (
// Equation(s):
// \RegWrite_EX~1_combout  = (instruction_D[31] & (instruction_D[30] $ ((instruction_D[28])))) # (!instruction_D[31] & (!instruction_D[30] & (instruction_D[28] $ (instruction_D[27]))))

	.dataa(instruction_D[31]),
	.datab(instruction_D[30]),
	.datac(instruction_D[28]),
	.datad(instruction_D[27]),
	.cin(gnd),
	.combout(\RegWrite_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \RegWrite_EX~1 .lut_mask = 16'h2938;
defparam \RegWrite_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N12
cycloneive_lcell_comb \RegWrite_EX~2 (
// Equation(s):
// \RegWrite_EX~2_combout  = (\RegWrite_EX~1_combout  & (((!\RegWrite_EX~0_combout  & !instruction_D[31])))) # (!\RegWrite_EX~1_combout  & (Decoder1 & ((instruction_D[31]))))

	.dataa(\CONTROL_UNIT|Decoder1~0_combout ),
	.datab(\RegWrite_EX~0_combout ),
	.datac(\RegWrite_EX~1_combout ),
	.datad(instruction_D[31]),
	.cin(gnd),
	.combout(\RegWrite_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \RegWrite_EX~2 .lut_mask = 16'h0A30;
defparam \RegWrite_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N14
cycloneive_lcell_comb \RegWrite_EX~3 (
// Equation(s):
// \RegWrite_EX~3_combout  = (\branch_or_jump~1_combout  & ((Equal31 & (Decoder0)) # (!Equal31 & ((!\RegWrite_EX~2_combout )))))

	.dataa(\branch_or_jump~1_combout ),
	.datab(\CONTROL_UNIT|Decoder0~1_combout ),
	.datac(\CONTROL_UNIT|Equal3~2_combout ),
	.datad(\RegWrite_EX~2_combout ),
	.cin(gnd),
	.combout(\RegWrite_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \RegWrite_EX~3 .lut_mask = 16'h808A;
defparam \RegWrite_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N20
cycloneive_lcell_comb \lui_EX~1 (
// Equation(s):
// \lui_EX~1_combout  = (\lui_EX~0_combout  & (instruction_D[29] & (instruction_D[28] & !instruction_D[31])))

	.dataa(\lui_EX~0_combout ),
	.datab(instruction_D[29]),
	.datac(instruction_D[28]),
	.datad(instruction_D[31]),
	.cin(gnd),
	.combout(\lui_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \lui_EX~1 .lut_mask = 16'h0080;
defparam \lui_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N25
dffeas \pc_plus_4_D[1] (
	.clk(CLK),
	.d(\pc_plus_4_D~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[1]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[1] .is_wysiwyg = "true";
defparam \pc_plus_4_D[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N12
cycloneive_lcell_comb \pc_plus_4_EX~0 (
// Equation(s):
// \pc_plus_4_EX~0_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[1] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_D[1]),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~0 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N0
cycloneive_lcell_comb \btbframes~2 (
// Equation(s):
// \btbframes~2_combout  = (\Mux29~1_combout  & (((\Mux30~1_combout  & !\always3~3_combout )) # (!\btbframes~0_combout ))) # (!\Mux29~1_combout  & (\Mux30~1_combout  & ((!\btbframes~0_combout ))))

	.dataa(\Mux29~1_combout ),
	.datab(\Mux30~1_combout ),
	.datac(\always3~3_combout ),
	.datad(\btbframes~0_combout ),
	.cin(gnd),
	.combout(\btbframes~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes~2 .lut_mask = 16'h08EE;
defparam \btbframes~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N14
cycloneive_lcell_comb \btbframes.frameblocks[3].curr_state[0]~1 (
// Equation(s):
// \btbframes.frameblocks[3].curr_state[0]~1_combout  = (!\branch_taken~0_combout  & (iwait & ((\Mux30~1_combout ) # (!\Mux29~1_combout ))))

	.dataa(\Mux29~1_combout ),
	.datab(\branch_taken~0_combout ),
	.datac(iwait),
	.datad(\Mux30~1_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].curr_state[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].curr_state[0]~1 .lut_mask = 16'h3010;
defparam \btbframes.frameblocks[3].curr_state[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N24
cycloneive_lcell_comb \btbframes.frameblocks[3].curr_state[0]~2 (
// Equation(s):
// \btbframes.frameblocks[3].curr_state[0]~2_combout  = (\nRST~input_o  & ((\btbframes.frameblocks[2].curr_state[0]~1_combout ) # ((\btbframes.frameblocks[3].curr_state[0]~1_combout  & \does_exist~18_combout ))))

	.dataa(\btbframes.frameblocks[2].curr_state[0]~1_combout ),
	.datab(nRST),
	.datac(\btbframes.frameblocks[3].curr_state[0]~1_combout ),
	.datad(\does_exist~18_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].curr_state[0]~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].curr_state[0]~2 .lut_mask = 16'hC888;
defparam \btbframes.frameblocks[3].curr_state[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N16
cycloneive_lcell_comb \btbframes.frameblocks[2].curr_state[0]~4 (
// Equation(s):
// \btbframes.frameblocks[2].curr_state[0]~4_combout  = (\Decoder0~0_combout  & ((\btbframes.frameblocks[3].curr_state[0]~2_combout  & (\btbframes~2_combout )) # (!\btbframes.frameblocks[3].curr_state[0]~2_combout  & ((\btbframes.frameblocks[2].curr_state 
// [0]))))) # (!\Decoder0~0_combout  & (((\btbframes.frameblocks[2].curr_state [0]))))

	.dataa(\Decoder0~0_combout ),
	.datab(\btbframes~2_combout ),
	.datac(\btbframes.frameblocks[2].curr_state [0]),
	.datad(\btbframes.frameblocks[3].curr_state[0]~2_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].curr_state[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].curr_state[0]~4 .lut_mask = 16'hD8F0;
defparam \btbframes.frameblocks[2].curr_state[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N10
cycloneive_lcell_comb \btbframes.frameblocks[1].curr_state[0]~3 (
// Equation(s):
// \btbframes.frameblocks[1].curr_state[0]~3_combout  = (\Decoder0~1_combout  & ((\btbframes.frameblocks[3].curr_state[0]~2_combout  & (\btbframes~2_combout )) # (!\btbframes.frameblocks[3].curr_state[0]~2_combout  & ((\btbframes.frameblocks[1].curr_state 
// [0]))))) # (!\Decoder0~1_combout  & (((\btbframes.frameblocks[1].curr_state [0]))))

	.dataa(\Decoder0~1_combout ),
	.datab(\btbframes~2_combout ),
	.datac(\btbframes.frameblocks[1].curr_state [0]),
	.datad(\btbframes.frameblocks[3].curr_state[0]~2_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].curr_state[0]~3_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].curr_state[0]~3 .lut_mask = 16'hD8F0;
defparam \btbframes.frameblocks[1].curr_state[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N20
cycloneive_lcell_comb \btbframes.frameblocks[0].curr_state[0]~3 (
// Equation(s):
// \btbframes.frameblocks[0].curr_state[0]~3_combout  = (\btbframes.frameblocks[0].curr_state[1]~1_combout  & (\btbframes~2_combout )) # (!\btbframes.frameblocks[0].curr_state[1]~1_combout  & ((\btbframes.frameblocks[0].curr_state [0])))

	.dataa(gnd),
	.datab(\btbframes~2_combout ),
	.datac(\btbframes.frameblocks[0].curr_state [0]),
	.datad(\btbframes.frameblocks[0].curr_state[1]~1_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].curr_state[0]~3_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].curr_state[0]~3 .lut_mask = 16'hCCF0;
defparam \btbframes.frameblocks[0].curr_state[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N12
cycloneive_lcell_comb \btbframes.frameblocks[3].curr_state[0]~3 (
// Equation(s):
// \btbframes.frameblocks[3].curr_state[0]~3_combout  = (\Decoder0~2_combout  & ((\btbframes.frameblocks[3].curr_state[0]~2_combout  & (\btbframes~2_combout )) # (!\btbframes.frameblocks[3].curr_state[0]~2_combout  & ((\btbframes.frameblocks[3].curr_state 
// [0]))))) # (!\Decoder0~2_combout  & (((\btbframes.frameblocks[3].curr_state [0]))))

	.dataa(\Decoder0~2_combout ),
	.datab(\btbframes~2_combout ),
	.datac(\btbframes.frameblocks[3].curr_state [0]),
	.datad(\btbframes.frameblocks[3].curr_state[0]~2_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].curr_state[0]~3_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].curr_state[0]~3 .lut_mask = 16'hD8F0;
defparam \btbframes.frameblocks[3].curr_state[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N23
dffeas \pc_plus_4_D[3] (
	.clk(CLK),
	.d(\pc_plus_4_D~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[3]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[3] .is_wysiwyg = "true";
defparam \pc_plus_4_D[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N13
dffeas \pc_plus_4_D[5] (
	.clk(CLK),
	.d(\pc_plus_4_D~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[5]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[5] .is_wysiwyg = "true";
defparam \pc_plus_4_D[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N27
dffeas \pc_plus_4_D[4] (
	.clk(CLK),
	.d(\pc_plus_4_D~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[4]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[4] .is_wysiwyg = "true";
defparam \pc_plus_4_D[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N23
dffeas \pc_plus_4_D[6] (
	.clk(CLK),
	.d(\pc_plus_4_D~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[6]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[6] .is_wysiwyg = "true";
defparam \pc_plus_4_D[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N5
dffeas \pc_plus_4_D[9] (
	.clk(CLK),
	.d(\pc_plus_4_D~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[9]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[9] .is_wysiwyg = "true";
defparam \pc_plus_4_D[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N27
dffeas \pc_plus_4_D[8] (
	.clk(CLK),
	.d(\pc_plus_4_D~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[8]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[8] .is_wysiwyg = "true";
defparam \pc_plus_4_D[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N20
cycloneive_lcell_comb \pc_plus_4_EX~9 (
// Equation(s):
// \pc_plus_4_EX~9_combout  = (pc_plus_4_D[8] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[8]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~9_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~9 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N13
dffeas \pc_plus_4_D[11] (
	.clk(CLK),
	.d(\pc_plus_4_D~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[11]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[11] .is_wysiwyg = "true";
defparam \pc_plus_4_D[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N13
dffeas \pc_plus_4_D[10] (
	.clk(CLK),
	.d(\pc_plus_4_D~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[10]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[10] .is_wysiwyg = "true";
defparam \pc_plus_4_D[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N11
dffeas \pc_plus_4_D[13] (
	.clk(CLK),
	.d(\pc_plus_4_D~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[13]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[13] .is_wysiwyg = "true";
defparam \pc_plus_4_D[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N3
dffeas \pc_plus_4_D[12] (
	.clk(CLK),
	.d(\pc_plus_4_D~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[12]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[12] .is_wysiwyg = "true";
defparam \pc_plus_4_D[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N14
cycloneive_lcell_comb \pc_plus_4_EX~13 (
// Equation(s):
// \pc_plus_4_EX~13_combout  = (pc_plus_4_D[12] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[12]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~13_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~13 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N11
dffeas \pc_plus_4_D[15] (
	.clk(CLK),
	.d(\pc_plus_4_D~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[15]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[15] .is_wysiwyg = "true";
defparam \pc_plus_4_D[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N2
cycloneive_lcell_comb \pc_plus_4_EX~14 (
// Equation(s):
// \pc_plus_4_EX~14_combout  = (pc_plus_4_D[15] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(pc_plus_4_D[15]),
	.datab(\branch_taken~0_combout ),
	.datac(\branch_or_jump~2_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~14_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~14 .lut_mask = 16'h8020;
defparam \pc_plus_4_EX~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N11
dffeas \pc_plus_4_D[14] (
	.clk(CLK),
	.d(\pc_plus_4_D~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[14]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[14] .is_wysiwyg = "true";
defparam \pc_plus_4_D[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N6
cycloneive_lcell_comb \pc_plus_4_EX~15 (
// Equation(s):
// \pc_plus_4_EX~15_combout  = (pc_plus_4_D[14] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[14]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~15_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~15 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N7
dffeas \pc_plus_4_D[16] (
	.clk(CLK),
	.d(\pc_plus_4_D~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[16]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[16] .is_wysiwyg = "true";
defparam \pc_plus_4_D[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N8
cycloneive_lcell_comb \pc_plus_4_EX~17 (
// Equation(s):
// \pc_plus_4_EX~17_combout  = (pc_plus_4_D[16] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_taken~0_combout ),
	.datab(pc_plus_4_D[16]),
	.datac(\predicted_M~q ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~17_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~17 .lut_mask = 16'h8400;
defparam \pc_plus_4_EX~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N7
dffeas \pc_plus_4_D[18] (
	.clk(CLK),
	.d(\pc_plus_4_D~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[18]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[18] .is_wysiwyg = "true";
defparam \pc_plus_4_D[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N16
cycloneive_lcell_comb \pc_plus_4_EX~19 (
// Equation(s):
// \pc_plus_4_EX~19_combout  = (pc_plus_4_D[18] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[18]),
	.datab(\predicted_M~q ),
	.datac(\branch_or_jump~2_combout ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~19_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~19 .lut_mask = 16'h8020;
defparam \pc_plus_4_EX~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N23
dffeas \pc_plus_4_D[21] (
	.clk(CLK),
	.d(\pc_plus_4_D~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[21]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[21] .is_wysiwyg = "true";
defparam \pc_plus_4_D[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N0
cycloneive_lcell_comb \pc_plus_4_EX~20 (
// Equation(s):
// \pc_plus_4_EX~20_combout  = (pc_plus_4_D[21] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(pc_plus_4_D[21]),
	.datab(\branch_taken~0_combout ),
	.datac(\branch_or_jump~2_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~20_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~20 .lut_mask = 16'h8020;
defparam \pc_plus_4_EX~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N5
dffeas \pc_plus_4_D[22] (
	.clk(CLK),
	.d(\pc_plus_4_D~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[22]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[22] .is_wysiwyg = "true";
defparam \pc_plus_4_D[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N22
cycloneive_lcell_comb \pc_plus_4_EX~23 (
// Equation(s):
// \pc_plus_4_EX~23_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[22] & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(\branch_taken~0_combout ),
	.datac(pc_plus_4_D[22]),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~23_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~23 .lut_mask = 16'h8020;
defparam \pc_plus_4_EX~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N31
dffeas \pc_plus_4_D[24] (
	.clk(CLK),
	.d(\pc_plus_4_D~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[24]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[24] .is_wysiwyg = "true";
defparam \pc_plus_4_D[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N27
dffeas \pc_plus_4_D[26] (
	.clk(CLK),
	.d(\pc_plus_4_D~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[26]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[26] .is_wysiwyg = "true";
defparam \pc_plus_4_D[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N27
dffeas \pc_plus_4_D[29] (
	.clk(CLK),
	.d(\pc_plus_4_D~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[29]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[29] .is_wysiwyg = "true";
defparam \pc_plus_4_D[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N24
cycloneive_lcell_comb \pc_plus_4_EX~28 (
// Equation(s):
// \pc_plus_4_EX~28_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[29] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(\predicted_M~q ),
	.datac(pc_plus_4_D[29]),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~28_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~28 .lut_mask = 16'h8020;
defparam \pc_plus_4_EX~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N3
dffeas \pc_plus_4_D[28] (
	.clk(CLK),
	.d(\pc_plus_4_D~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[28]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[28] .is_wysiwyg = "true";
defparam \pc_plus_4_D[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N30
cycloneive_lcell_comb \pc_plus_4_EX~29 (
// Equation(s):
// \pc_plus_4_EX~29_combout  = (pc_plus_4_D[28] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(pc_plus_4_D[28]),
	.datac(\branch_taken~0_combout ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~29_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~29 .lut_mask = 16'h8400;
defparam \pc_plus_4_EX~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N11
dffeas \pc_plus_4_D[31] (
	.clk(CLK),
	.d(\pc_plus_4_D~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[31]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[31] .is_wysiwyg = "true";
defparam \pc_plus_4_D[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N10
cycloneive_lcell_comb \predicted_D~0 (
// Equation(s):
// \predicted_D~0_combout  = (\branch_or_jump~1_combout  & (iwait & predicted))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(iwait),
	.datad(\BTB|predicted~18_combout ),
	.cin(gnd),
	.combout(\predicted_D~0_combout ),
	.cout());
// synopsys translate_off
defparam \predicted_D~0 .lut_mask = 16'hA000;
defparam \predicted_D~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N24
cycloneive_lcell_comb \pc_plus_4_D~0 (
// Equation(s):
// \pc_plus_4_D~0_combout  = (pc_out_1 & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(pc_out_1),
	.cin(gnd),
	.combout(\pc_plus_4_D~0_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~0 .lut_mask = 16'hF300;
defparam \pc_plus_4_D~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N22
cycloneive_lcell_comb \pc_plus_4_D~2 (
// Equation(s):
// \pc_plus_4_D~2_combout  = (\pc_plus_4[3]~2_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(\pc_plus_4[3]~2_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\pc_plus_4_D~2_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~2 .lut_mask = 16'hF050;
defparam \pc_plus_4_D~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N12
cycloneive_lcell_comb \pc_plus_4_D~4 (
// Equation(s):
// \pc_plus_4_D~4_combout  = (\pc_plus_4[5]~6_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\pc_plus_4[5]~6_combout ),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_plus_4_D~4_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~4 .lut_mask = 16'hA2A2;
defparam \pc_plus_4_D~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N26
cycloneive_lcell_comb \pc_plus_4_D~5 (
// Equation(s):
// \pc_plus_4_D~5_combout  = (\pc_plus_4[4]~4_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\pc_plus_4[4]~4_combout ),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\pc_plus_4_D~5_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~5 .lut_mask = 16'hAA0A;
defparam \pc_plus_4_D~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N22
cycloneive_lcell_comb \pc_plus_4_D~7 (
// Equation(s):
// \pc_plus_4_D~7_combout  = (\pc_plus_4[6]~8_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(\pc_plus_4[6]~8_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\pc_plus_4_D~7_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~7 .lut_mask = 16'hF030;
defparam \pc_plus_4_D~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N4
cycloneive_lcell_comb \pc_plus_4_D~8 (
// Equation(s):
// \pc_plus_4_D~8_combout  = (\pc_plus_4[9]~14_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(iwait),
	.datab(\branch_or_jump~1_combout ),
	.datac(gnd),
	.datad(\pc_plus_4[9]~14_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~8_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~8 .lut_mask = 16'hBB00;
defparam \pc_plus_4_D~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N26
cycloneive_lcell_comb \pc_plus_4_D~9 (
// Equation(s):
// \pc_plus_4_D~9_combout  = (\pc_plus_4[8]~12_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(\pc_plus_4[8]~12_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\pc_plus_4_D~9_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~9 .lut_mask = 16'hF030;
defparam \pc_plus_4_D~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N12
cycloneive_lcell_comb \pc_plus_4_D~10 (
// Equation(s):
// \pc_plus_4_D~10_combout  = (\pc_plus_4[11]~18_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(iwait),
	.datad(\pc_plus_4[11]~18_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~10_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~10 .lut_mask = 16'hF500;
defparam \pc_plus_4_D~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N12
cycloneive_lcell_comb \pc_plus_4_D~11 (
// Equation(s):
// \pc_plus_4_D~11_combout  = (\pc_plus_4[10]~16_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(gnd),
	.datab(iwait),
	.datac(\branch_or_jump~1_combout ),
	.datad(\pc_plus_4[10]~16_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~11_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~11 .lut_mask = 16'hCF00;
defparam \pc_plus_4_D~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N10
cycloneive_lcell_comb \pc_plus_4_D~12 (
// Equation(s):
// \pc_plus_4_D~12_combout  = (\pc_plus_4[13]~22_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(gnd),
	.datab(iwait),
	.datac(\pc_plus_4[13]~22_combout ),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~12_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~12 .lut_mask = 16'hC0F0;
defparam \pc_plus_4_D~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N2
cycloneive_lcell_comb \pc_plus_4_D~13 (
// Equation(s):
// \pc_plus_4_D~13_combout  = (\pc_plus_4[12]~20_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(gnd),
	.datab(iwait),
	.datac(\pc_plus_4[12]~20_combout ),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~13_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~13 .lut_mask = 16'hC0F0;
defparam \pc_plus_4_D~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N10
cycloneive_lcell_comb \pc_plus_4_D~14 (
// Equation(s):
// \pc_plus_4_D~14_combout  = (\pc_plus_4[15]~26_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(iwait),
	.datab(\pc_plus_4[15]~26_combout ),
	.datac(gnd),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~14_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~14 .lut_mask = 16'h88CC;
defparam \pc_plus_4_D~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N10
cycloneive_lcell_comb \pc_plus_4_D~15 (
// Equation(s):
// \pc_plus_4_D~15_combout  = (\pc_plus_4[14]~24_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(iwait),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\pc_plus_4[14]~24_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~15_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~15 .lut_mask = 16'hAF00;
defparam \pc_plus_4_D~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N6
cycloneive_lcell_comb \pc_plus_4_D~17 (
// Equation(s):
// \pc_plus_4_D~17_combout  = (\pc_plus_4[16]~28_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\pc_plus_4[16]~28_combout ),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_plus_4_D~17_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~17 .lut_mask = 16'hA2A2;
defparam \pc_plus_4_D~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N6
cycloneive_lcell_comb \pc_plus_4_D~19 (
// Equation(s):
// \pc_plus_4_D~19_combout  = (\pc_plus_4[18]~32_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\pc_plus_4[18]~32_combout ),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_plus_4_D~19_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~19 .lut_mask = 16'hA2A2;
defparam \pc_plus_4_D~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N22
cycloneive_lcell_comb \pc_plus_4_D~20 (
// Equation(s):
// \pc_plus_4_D~20_combout  = (\pc_plus_4[21]~38_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(iwait),
	.datab(gnd),
	.datac(\pc_plus_4[21]~38_combout ),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~20_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~20 .lut_mask = 16'hA0F0;
defparam \pc_plus_4_D~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N4
cycloneive_lcell_comb \pc_plus_4_D~23 (
// Equation(s):
// \pc_plus_4_D~23_combout  = (\pc_plus_4[22]~40_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\pc_plus_4[22]~40_combout ),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_plus_4_D~23_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~23 .lut_mask = 16'hA2A2;
defparam \pc_plus_4_D~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N30
cycloneive_lcell_comb \pc_plus_4_D~25 (
// Equation(s):
// \pc_plus_4_D~25_combout  = (\pc_plus_4[24]~44_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(\pc_plus_4[24]~44_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\pc_plus_4_D~25_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~25 .lut_mask = 16'hF050;
defparam \pc_plus_4_D~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N26
cycloneive_lcell_comb \pc_plus_4_D~27 (
// Equation(s):
// \pc_plus_4_D~27_combout  = (\pc_plus_4[26]~48_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(iwait),
	.datab(\branch_or_jump~1_combout ),
	.datac(gnd),
	.datad(\pc_plus_4[26]~48_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~27_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~27 .lut_mask = 16'hBB00;
defparam \pc_plus_4_D~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N26
cycloneive_lcell_comb \pc_plus_4_D~28 (
// Equation(s):
// \pc_plus_4_D~28_combout  = (\pc_plus_4[29]~54_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(\pc_plus_4[29]~54_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~28_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~28 .lut_mask = 16'hF300;
defparam \pc_plus_4_D~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N2
cycloneive_lcell_comb \pc_plus_4_D~29 (
// Equation(s):
// \pc_plus_4_D~29_combout  = (\pc_plus_4[28]~52_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\branch_or_jump~1_combout ),
	.datab(\pc_plus_4[28]~52_combout ),
	.datac(iwait),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_plus_4_D~29_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~29 .lut_mask = 16'hC4C4;
defparam \pc_plus_4_D~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N10
cycloneive_lcell_comb \pc_plus_4_D~30 (
// Equation(s):
// \pc_plus_4_D~30_combout  = (\pc_plus_4[31]~58_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(\pc_plus_4[31]~58_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\pc_plus_4_D~30_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~30 .lut_mask = 16'hF050;
defparam \pc_plus_4_D~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N0
cycloneive_lcell_comb \portB~112 (
// Equation(s):
// \portB~112_combout  = (\portB~14_combout  & (!\lui_M~q  & ((porto_M_13)))) # (!\portB~14_combout  & (((\wdat_WB[13]~39_combout ))))

	.dataa(\lui_M~q ),
	.datab(\wdat_WB[13]~39_combout ),
	.datac(porto_M_13),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~112_combout ),
	.cout());
// synopsys translate_off
defparam \portB~112 .lut_mask = 16'h50CC;
defparam \portB~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N10
cycloneive_lcell_comb \portB~113 (
// Equation(s):
// \portB~113_combout  = (\portB~14_combout  & (!\lui_M~q  & ((porto_M_12)))) # (!\portB~14_combout  & (((\wdat_WB[12]~41_combout ))))

	.dataa(\lui_M~q ),
	.datab(\wdat_WB[12]~41_combout ),
	.datac(porto_M_12),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~113_combout ),
	.cout());
// synopsys translate_off
defparam \portB~113 .lut_mask = 16'h50CC;
defparam \portB~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N8
cycloneive_lcell_comb \portB~114 (
// Equation(s):
// \portB~114_combout  = (\portB~14_combout  & (!\lui_M~q  & (porto_M_7))) # (!\portB~14_combout  & (((\wdat_WB[7]~51_combout ))))

	.dataa(\lui_M~q ),
	.datab(porto_M_7),
	.datac(\wdat_WB[7]~51_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~114_combout ),
	.cout());
// synopsys translate_off
defparam \portB~114 .lut_mask = 16'h44F0;
defparam \portB~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N10
cycloneive_lcell_comb \portB~116 (
// Equation(s):
// \portB~116_combout  = (\Equal2~0_combout  & (porto_M_5 & (!\lui_M~q ))) # (!\Equal2~0_combout  & (((\portB~86_combout ))))

	.dataa(porto_M_5),
	.datab(\lui_M~q ),
	.datac(\Equal2~0_combout ),
	.datad(\portB~86_combout ),
	.cin(gnd),
	.combout(\portB~116_combout ),
	.cout());
// synopsys translate_off
defparam \portB~116 .lut_mask = 16'h2F20;
defparam \portB~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N18
cycloneive_lcell_comb \portA~70 (
// Equation(s):
// \portA~70_combout  = (fuifforward_A_01 & (((porto_M_8 & !\lui_M~q )))) # (!fuifforward_A_01 & (rdata1_EX[8]))

	.dataa(rdata1_EX[8]),
	.datab(porto_M_8),
	.datac(\lui_M~q ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~70_combout ),
	.cout());
// synopsys translate_off
defparam \portA~70 .lut_mask = 16'h0CAA;
defparam \portA~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N18
cycloneive_lcell_comb \portA~71 (
// Equation(s):
// \portA~71_combout  = (fuifforward_A_01 & (porto_M_10 & (!\lui_M~q ))) # (!fuifforward_A_01 & (((rdata1_EX[10]))))

	.dataa(porto_M_10),
	.datab(\lui_M~q ),
	.datac(rdata1_EX[10]),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~71_combout ),
	.cout());
// synopsys translate_off
defparam \portA~71 .lut_mask = 16'h22F0;
defparam \portA~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N30
cycloneive_lcell_comb \portA~72 (
// Equation(s):
// \portA~72_combout  = (fuifforward_A_01 & (((porto_M_9 & !\lui_M~q )))) # (!fuifforward_A_01 & (rdata1_EX[9]))

	.dataa(rdata1_EX[9]),
	.datab(porto_M_9),
	.datac(\lui_M~q ),
	.datad(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.cin(gnd),
	.combout(\portA~72_combout ),
	.cout());
// synopsys translate_off
defparam \portA~72 .lut_mask = 16'h0CAA;
defparam \portA~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N16
cycloneive_lcell_comb \comb~3 (
// Equation(s):
// \comb~3_combout  = (!dREN_M1 & (!dWEN_M1 & (always1 & !Decoder11)))

	.dataa(dREN_M1),
	.datab(dWEN_M1),
	.datac(always1),
	.datad(\CONTROL_UNIT|Decoder1~1_combout ),
	.cin(gnd),
	.combout(\comb~3_combout ),
	.cout());
// synopsys translate_off
defparam \comb~3 .lut_mask = 16'h0010;
defparam \comb~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N2
cycloneive_lcell_comb \btbframes.frameblocks[2].tag[27]~3 (
// Equation(s):
// \btbframes.frameblocks[2].tag[27]~3_combout  = (\nRST~input_o  & ((\beq_M~q ) # (\bne_M~q )))

	.dataa(gnd),
	.datab(\beq_M~q ),
	.datac(\bne_M~q ),
	.datad(nRST),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].tag[27]~3_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[27]~3 .lut_mask = 16'hFC00;
defparam \btbframes.frameblocks[2].tag[27]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N20
cycloneive_lcell_comb \btbframes.frameblocks[0].tag[27]~3 (
// Equation(s):
// \btbframes.frameblocks[0].tag[27]~3_combout  = (!\Add2~2_combout  & (\nRST~input_o  & ((\beq_M~q ) # (\bne_M~q ))))

	.dataa(\Add2~2_combout ),
	.datab(\beq_M~q ),
	.datac(\bne_M~q ),
	.datad(nRST),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].tag[27]~3_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[27]~3 .lut_mask = 16'h5400;
defparam \btbframes.frameblocks[0].tag[27]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N16
cycloneive_lcell_comb \always3~3 (
// Equation(s):
// \always3~3_combout  = (iwait & (!\does_exist~18_combout  & ((\bne_M~q ) # (\beq_M~q ))))

	.dataa(\bne_M~q ),
	.datab(\beq_M~q ),
	.datac(iwait),
	.datad(\does_exist~18_combout ),
	.cin(gnd),
	.combout(\always3~3_combout ),
	.cout());
// synopsys translate_off
defparam \always3~3 .lut_mask = 16'h00E0;
defparam \always3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N2
cycloneive_lcell_comb \btbframes.frameblocks[2].valid~2 (
// Equation(s):
// \btbframes.frameblocks[2].valid~2_combout  = (\btbframes.frameblocks[2].valid~q ) # ((\Add2~2_combout  & (\always3~3_combout  & !\Add2~0_combout )))

	.dataa(\Add2~2_combout ),
	.datab(\always3~3_combout ),
	.datac(\btbframes.frameblocks[2].valid~q ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].valid~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].valid~2 .lut_mask = 16'hF0F8;
defparam \btbframes.frameblocks[2].valid~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N20
cycloneive_lcell_comb \btbframes.frameblocks[1].valid~2 (
// Equation(s):
// \btbframes.frameblocks[1].valid~2_combout  = (\btbframes.frameblocks[1].valid~q ) # ((!\Add2~2_combout  & (\always3~3_combout  & \Add2~0_combout )))

	.dataa(\Add2~2_combout ),
	.datab(\always3~3_combout ),
	.datac(\btbframes.frameblocks[1].valid~q ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].valid~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].valid~2 .lut_mask = 16'hF4F0;
defparam \btbframes.frameblocks[1].valid~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N14
cycloneive_lcell_comb \btbframes.frameblocks[3].valid~2 (
// Equation(s):
// \btbframes.frameblocks[3].valid~2_combout  = (\btbframes.frameblocks[3].valid~q ) # ((\Add2~2_combout  & (\always3~3_combout  & \Add2~0_combout )))

	.dataa(\Add2~2_combout ),
	.datab(\always3~3_combout ),
	.datac(\btbframes.frameblocks[3].valid~q ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].valid~2_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].valid~2 .lut_mask = 16'hF8F0;
defparam \btbframes.frameblocks[3].valid~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N20
cycloneive_lcell_comb \jal_EX~2 (
// Equation(s):
// \jal_EX~2_combout  = (!instruction_D[31] & (!instruction_D[29] & (\lui_EX~0_combout  & !instruction_D[28])))

	.dataa(instruction_D[31]),
	.datab(instruction_D[29]),
	.datac(\lui_EX~0_combout ),
	.datad(instruction_D[28]),
	.cin(gnd),
	.combout(\jal_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \jal_EX~2 .lut_mask = 16'h0010;
defparam \jal_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N28
cycloneive_lcell_comb \instruction_D~70 (
// Equation(s):
// \instruction_D~70_combout  = (\branch_or_jump~1_combout  & (ramiframload_16 & iwait))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(\dpif.dmemload [16]),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~70_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~70 .lut_mask = 16'hC000;
defparam \instruction_D~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N0
cycloneive_lcell_comb \instruction_D~71 (
// Equation(s):
// \instruction_D~71_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_17))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(iwait),
	.datad(\dpif.dmemload [17]),
	.cin(gnd),
	.combout(\instruction_D~71_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~71 .lut_mask = 16'hA000;
defparam \instruction_D~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N6
cycloneive_lcell_comb \instruction_D~72 (
// Equation(s):
// \instruction_D~72_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_18))

	.dataa(\branch_or_jump~1_combout ),
	.datab(iwait),
	.datac(ramiframload_18),
	.datad(gnd),
	.cin(gnd),
	.combout(\instruction_D~72_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~72 .lut_mask = 16'h8080;
defparam \instruction_D~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N30
cycloneive_lcell_comb \instruction_D~73 (
// Equation(s):
// \instruction_D~73_combout  = (\branch_or_jump~1_combout  & (ramiframload_19 & iwait))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(ramiframload_19),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~73_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~73 .lut_mask = 16'hC000;
defparam \instruction_D~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N8
cycloneive_lcell_comb \instruction_D~75 (
// Equation(s):
// \instruction_D~75_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_22))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(ramiframload_22),
	.cin(gnd),
	.combout(\instruction_D~75_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~75 .lut_mask = 16'hC000;
defparam \instruction_D~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N8
cycloneive_lcell_comb \instruction_D~77 (
// Equation(s):
// \instruction_D~77_combout  = (\branch_or_jump~1_combout  & (ramiframload_24 & iwait))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(ramiframload_24),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~77_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~77 .lut_mask = 16'hC000;
defparam \instruction_D~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N14
cycloneive_lcell_comb \instruction_D~78 (
// Equation(s):
// \instruction_D~78_combout  = (iwait & (ramiframload_23 & \branch_or_jump~1_combout ))

	.dataa(iwait),
	.datab(\dpif.dmemload [23]),
	.datac(gnd),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\instruction_D~78_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~78 .lut_mask = 16'h8800;
defparam \instruction_D~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N12
cycloneive_lcell_comb \instruction_D~79 (
// Equation(s):
// \instruction_D~79_combout  = (ramiframload_25 & (iwait & \branch_or_jump~1_combout ))

	.dataa(gnd),
	.datab(\dpif.dmemload [25]),
	.datac(iwait),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\instruction_D~79_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~79 .lut_mask = 16'hC000;
defparam \instruction_D~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N4
cycloneive_lcell_comb \instruction_D~92 (
// Equation(s):
// \instruction_D~92_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_11))

	.dataa(\branch_or_jump~1_combout ),
	.datab(iwait),
	.datac(gnd),
	.datad(\dpif.dmemload [11]),
	.cin(gnd),
	.combout(\instruction_D~92_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~92 .lut_mask = 16'h8800;
defparam \instruction_D~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N8
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[3]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[3]~feeder_combout  = \pc_when_branch[3]~2_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[3]~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[3]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[1].jump_add[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N24
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[3]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[3]~feeder_combout  = \pc_when_branch[3]~2_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[3]~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[3]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].jump_add[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N28
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[4]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[4]~feeder_combout  = \pc_when_branch[4]~4_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[4]~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[4]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[1].jump_add[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N24
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[6]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[6]~feeder_combout  = \pc_when_branch[6]~8_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[6]~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[6]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].jump_add[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N10
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[7]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[7]~feeder_combout  = \pc_when_branch[7]~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[7]~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[7]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[1].jump_add[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N26
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[8]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[8]~feeder_combout  = \pc_when_branch[8]~12_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[8]~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[8]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].jump_add[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N30
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[10]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[10]~feeder_combout  = \pc_when_branch[10]~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[10]~16_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[10]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].jump_add[10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N16
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[10]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[10]~feeder_combout  = \pc_when_branch[10]~16_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[10]~16_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[10]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[1].jump_add[10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N0
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[11]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[11]~feeder_combout  = \pc_when_branch[11]~18_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[11]~18_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[11]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[2].jump_add[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N28
cycloneive_lcell_comb \btbframes.frameblocks[0].jump_add[11]~feeder (
// Equation(s):
// \btbframes.frameblocks[0].jump_add[11]~feeder_combout  = \pc_when_branch[11]~18_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[11]~18_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].jump_add[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[11]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[0].jump_add[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N24
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[12]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[12]~feeder_combout  = \pc_when_branch[12]~20_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[12]~20_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[12]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[1].jump_add[12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N26
cycloneive_lcell_comb \btbframes.frameblocks[0].jump_add[13]~feeder (
// Equation(s):
// \btbframes.frameblocks[0].jump_add[13]~feeder_combout  = \pc_when_branch[13]~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[13]~22_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].jump_add[13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[13]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[0].jump_add[13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N20
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[13]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[13]~feeder_combout  = \pc_when_branch[13]~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[13]~22_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[13]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].jump_add[13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N24
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[14]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[14]~feeder_combout  = \pc_when_branch[14]~24_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[14]~24_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[14]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[1].jump_add[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N16
cycloneive_lcell_comb \btbframes.frameblocks[0].jump_add[14]~feeder (
// Equation(s):
// \btbframes.frameblocks[0].jump_add[14]~feeder_combout  = \pc_when_branch[14]~24_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[14]~24_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].jump_add[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[14]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[0].jump_add[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N20
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[15]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[15]~feeder_combout  = \pc_when_branch[15]~26_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[15]~26_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[15]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[1].jump_add[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N8
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[16]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[16]~feeder_combout  = \pc_when_branch[16]~28_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[16]~28_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[16]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].jump_add[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N10
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[16]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[16]~feeder_combout  = \pc_when_branch[16]~28_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[16]~28_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[16]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[1].jump_add[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N14
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[18]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[18]~feeder_combout  = \pc_when_branch[18]~32_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[18]~32_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[18]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[2].jump_add[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N18
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[19]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[19]~feeder_combout  = \pc_when_branch[19]~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[19]~34_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[19]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].jump_add[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N2
cycloneive_lcell_comb \btbframes.frameblocks[0].jump_add[20]~feeder (
// Equation(s):
// \btbframes.frameblocks[0].jump_add[20]~feeder_combout  = \pc_when_branch[20]~36_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[20]~36_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].jump_add[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].jump_add[20]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[0].jump_add[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N4
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[21]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[21]~feeder_combout  = \pc_when_branch[21]~38_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[21]~38_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[21]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[1].jump_add[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N14
cycloneive_lcell_comb \btbframes.frameblocks[3].jump_add[21]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].jump_add[21]~feeder_combout  = \pc_when_branch[21]~38_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[21]~38_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].jump_add[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[21]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[3].jump_add[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N0
cycloneive_lcell_comb \btbframes.frameblocks[3].jump_add[23]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].jump_add[23]~feeder_combout  = \pc_when_branch[23]~42_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[23]~42_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].jump_add[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[23]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[3].jump_add[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N20
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[23]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[23]~feeder_combout  = \pc_when_branch[23]~42_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[23]~42_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[23]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[1].jump_add[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N16
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[24]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[24]~feeder_combout  = \pc_when_branch[24]~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[24]~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[24]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].jump_add[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N0
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[26]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[26]~feeder_combout  = \pc_when_branch[26]~48_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[26]~48_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[26]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].jump_add[26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N28
cycloneive_lcell_comb \btbframes.frameblocks[3].jump_add[26]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].jump_add[26]~feeder_combout  = \pc_when_branch[26]~48_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\pc_when_branch[26]~48_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].jump_add[26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].jump_add[26]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[3].jump_add[26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N30
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[28]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[28]~feeder_combout  = \pc_when_branch[28]~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[28]~52_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[28]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[1].jump_add[28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N16
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[28]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[28]~feeder_combout  = \pc_when_branch[28]~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[28]~52_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[28]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[2].jump_add[28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N12
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[30]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[30]~feeder_combout  = \pc_when_branch[30]~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[30]~56_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[30]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[2].jump_add[30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N14
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[31]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[31]~feeder_combout  = \pc_when_branch[31]~58_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\pc_when_branch[31]~58_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[31]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[2].jump_add[31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N6
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[0]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[0]~feeder_combout  = \Add2~4_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[0]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[3].tag[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N0
cycloneive_lcell_comb \btbframes.frameblocks[0].tag[1]~feeder (
// Equation(s):
// \btbframes.frameblocks[0].tag[1]~feeder_combout  = \Add2~6_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].tag[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[1]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[0].tag[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N20
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[2]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[2]~feeder_combout  = \Add2~8_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[2]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[3].tag[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N4
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[3]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[3]~feeder_combout  = \Add2~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add2~10_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[3]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[3].tag[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N2
cycloneive_lcell_comb \btbframes.frameblocks[0].tag[3]~feeder (
// Equation(s):
// \btbframes.frameblocks[0].tag[3]~feeder_combout  = \Add2~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].tag[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[3]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[0].tag[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N18
cycloneive_lcell_comb \btbframes.frameblocks[2].tag[5]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].tag[5]~feeder_combout  = \Add2~14_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].tag[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[5]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].tag[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N16
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[8]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[8]~feeder_combout  = \Add2~20_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~20_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[8]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[3].tag[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N16
cycloneive_lcell_comb \btbframes.frameblocks[1].tag[9]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].tag[9]~feeder_combout  = \Add2~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add2~22_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].tag[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[9]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[1].tag[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N10
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[9]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[9]~feeder_combout  = \Add2~22_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add2~22_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[9]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[3].tag[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N2
cycloneive_lcell_comb \btbframes.frameblocks[1].tag[15]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].tag[15]~feeder_combout  = \Add2~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add2~34_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].tag[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[15]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[1].tag[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N26
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[15]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[15]~feeder_combout  = \Add2~34_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~34_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[15]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[3].tag[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N4
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[16]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[16]~feeder_combout  = \Add2~36_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~36_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[16]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[3].tag[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N16
cycloneive_lcell_comb \btbframes.frameblocks[2].tag[16]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].tag[16]~feeder_combout  = \Add2~36_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add2~36_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].tag[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[16]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[2].tag[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N28
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[18]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[18]~feeder_combout  = \Add2~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~40_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[18]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[3].tag[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N0
cycloneive_lcell_comb \btbframes.frameblocks[1].tag[18]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].tag[18]~feeder_combout  = \Add2~40_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~40_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].tag[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[18]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[1].tag[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N20
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[20]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[20]~feeder_combout  = \Add2~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[20]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[3].tag[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N30
cycloneive_lcell_comb \btbframes.frameblocks[2].tag[20]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].tag[20]~feeder_combout  = \Add2~44_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~44_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].tag[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[20]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].tag[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N2
cycloneive_lcell_comb \btbframes.frameblocks[0].tag[21]~feeder (
// Equation(s):
// \btbframes.frameblocks[0].tag[21]~feeder_combout  = \Add2~46_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~46_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].tag[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[21]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[0].tag[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N2
cycloneive_lcell_comb \btbframes.frameblocks[2].tag[22]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].tag[22]~feeder_combout  = \Add2~48_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add2~48_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].tag[22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[22]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[2].tag[22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N22
cycloneive_lcell_comb \btbframes.frameblocks[1].tag[23]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].tag[23]~feeder_combout  = \Add2~50_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~50_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].tag[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].tag[23]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[1].tag[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N30
cycloneive_lcell_comb \btbframes.frameblocks[0].tag[24]~feeder (
// Equation(s):
// \btbframes.frameblocks[0].tag[24]~feeder_combout  = \Add2~52_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~52_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[0].tag[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[0].tag[24]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[0].tag[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N26
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[26]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[26]~feeder_combout  = \Add2~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~56_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[26]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[3].tag[26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N0
cycloneive_lcell_comb \btbframes.frameblocks[2].tag[26]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].tag[26]~feeder_combout  = \Add2~56_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add2~56_combout ),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].tag[26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].tag[26]~feeder .lut_mask = 16'hFF00;
defparam \btbframes.frameblocks[2].tag[26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N28
cycloneive_lcell_comb \btbframes.frameblocks[3].tag[27]~feeder (
// Equation(s):
// \btbframes.frameblocks[3].tag[27]~feeder_combout  = \Add2~58_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add2~58_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[3].tag[27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[3].tag[27]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[3].tag[27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N4
cycloneive_lcell_comb \dmemload_WB[4]~feeder (
// Equation(s):
// \dmemload_WB[4]~feeder_combout  = ramiframload_4

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_4),
	.cin(gnd),
	.combout(\dmemload_WB[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \dmemload_WB[4]~feeder .lut_mask = 16'hFF00;
defparam \dmemload_WB[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N0
cycloneive_lcell_comb \dmemload_WB[15]~feeder (
// Equation(s):
// \dmemload_WB[15]~feeder_combout  = ramiframload_15

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_15),
	.cin(gnd),
	.combout(\dmemload_WB[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \dmemload_WB[15]~feeder .lut_mask = 16'hFF00;
defparam \dmemload_WB[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N30
cycloneive_lcell_comb \dmemload_WB[18]~feeder (
// Equation(s):
// \dmemload_WB[18]~feeder_combout  = ramiframload_18

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_18),
	.cin(gnd),
	.combout(\dmemload_WB[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \dmemload_WB[18]~feeder .lut_mask = 16'hFF00;
defparam \dmemload_WB[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N22
cycloneive_lcell_comb \dmemload_WB[19]~feeder (
// Equation(s):
// \dmemload_WB[19]~feeder_combout  = ramiframload_19

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_19),
	.cin(gnd),
	.combout(\dmemload_WB[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \dmemload_WB[19]~feeder .lut_mask = 16'hFF00;
defparam \dmemload_WB[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N16
cycloneive_lcell_comb \btbframes.frameblocks[2].jump_add[1]~feeder (
// Equation(s):
// \btbframes.frameblocks[2].jump_add[1]~feeder_combout  = pc_plus_4_M[1]

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_plus_4_M[1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[2].jump_add[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[2].jump_add[1]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[2].jump_add[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N12
cycloneive_lcell_comb \btbframes.frameblocks[1].jump_add[0]~feeder (
// Equation(s):
// \btbframes.frameblocks[1].jump_add[0]~feeder_combout  = pc_plus_4_M[0]

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_plus_4_M[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\btbframes.frameblocks[1].jump_add[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \btbframes.frameblocks[1].jump_add[0]~feeder .lut_mask = 16'hF0F0;
defparam \btbframes.frameblocks[1].jump_add[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N12
cycloneive_lcell_comb \pc_plus_4_WB[18]~feeder (
// Equation(s):
// \pc_plus_4_WB[18]~feeder_combout  = pc_plus_4_M[18]

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pc_plus_4_M[18]),
	.cin(gnd),
	.combout(\pc_plus_4_WB[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_WB[18]~feeder .lut_mask = 16'hFF00;
defparam \pc_plus_4_WB[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N5
dffeas \rdata2_M[0] (
	.clk(CLK),
	.d(\rdata2_M~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_0),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[0] .is_wysiwyg = "true";
defparam \rdata2_M[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N9
dffeas \rdata2_M[1] (
	.clk(CLK),
	.d(\rdata2_M~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_1),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[1] .is_wysiwyg = "true";
defparam \rdata2_M[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N25
dffeas \rdata2_M[2] (
	.clk(CLK),
	.d(\rdata2_M~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_2),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[2] .is_wysiwyg = "true";
defparam \rdata2_M[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N1
dffeas \rdata2_M[3] (
	.clk(CLK),
	.d(\rdata2_M~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_3),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[3] .is_wysiwyg = "true";
defparam \rdata2_M[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N21
dffeas \rdata2_M[4] (
	.clk(CLK),
	.d(\rdata2_M~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_4),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[4] .is_wysiwyg = "true";
defparam \rdata2_M[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N1
dffeas \rdata2_M[5] (
	.clk(CLK),
	.d(\rdata2_M~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_5),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[5] .is_wysiwyg = "true";
defparam \rdata2_M[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N11
dffeas \rdata2_M[6] (
	.clk(CLK),
	.d(\rdata2_M~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_6),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[6] .is_wysiwyg = "true";
defparam \rdata2_M[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N15
dffeas \rdata2_M[7] (
	.clk(CLK),
	.d(\rdata2_M~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_7),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[7] .is_wysiwyg = "true";
defparam \rdata2_M[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N13
dffeas \rdata2_M[8] (
	.clk(CLK),
	.d(\rdata2_M~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_8),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[8] .is_wysiwyg = "true";
defparam \rdata2_M[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N21
dffeas \rdata2_M[9] (
	.clk(CLK),
	.d(\rdata2_M~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_9),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[9] .is_wysiwyg = "true";
defparam \rdata2_M[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N3
dffeas \rdata2_M[10] (
	.clk(CLK),
	.d(\rdata2_M~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_10),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[10] .is_wysiwyg = "true";
defparam \rdata2_M[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N7
dffeas \rdata2_M[11] (
	.clk(CLK),
	.d(\rdata2_M~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_11),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[11] .is_wysiwyg = "true";
defparam \rdata2_M[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N23
dffeas \rdata2_M[12] (
	.clk(CLK),
	.d(\rdata2_M~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_12),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[12] .is_wysiwyg = "true";
defparam \rdata2_M[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N9
dffeas \rdata2_M[13] (
	.clk(CLK),
	.d(\rdata2_M~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_13),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[13] .is_wysiwyg = "true";
defparam \rdata2_M[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N25
dffeas \rdata2_M[14] (
	.clk(CLK),
	.d(\rdata2_M~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_14),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[14] .is_wysiwyg = "true";
defparam \rdata2_M[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N21
dffeas \rdata2_M[15] (
	.clk(CLK),
	.d(\rdata2_M~33_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_15),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[15] .is_wysiwyg = "true";
defparam \rdata2_M[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N11
dffeas \rdata2_M[16] (
	.clk(CLK),
	.d(\rdata2_M~35_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_16),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[16] .is_wysiwyg = "true";
defparam \rdata2_M[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N25
dffeas \rdata2_M[17] (
	.clk(CLK),
	.d(\rdata2_M~37_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_17),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[17] .is_wysiwyg = "true";
defparam \rdata2_M[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N17
dffeas \rdata2_M[18] (
	.clk(CLK),
	.d(\rdata2_M~39_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_18),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[18] .is_wysiwyg = "true";
defparam \rdata2_M[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N3
dffeas \rdata2_M[19] (
	.clk(CLK),
	.d(\rdata2_M~41_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_19),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[19] .is_wysiwyg = "true";
defparam \rdata2_M[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N1
dffeas \rdata2_M[20] (
	.clk(CLK),
	.d(\rdata2_M~43_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_20),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[20] .is_wysiwyg = "true";
defparam \rdata2_M[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N11
dffeas \rdata2_M[21] (
	.clk(CLK),
	.d(\rdata2_M~45_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_21),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[21] .is_wysiwyg = "true";
defparam \rdata2_M[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N11
dffeas \rdata2_M[22] (
	.clk(CLK),
	.d(\rdata2_M~47_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_22),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[22] .is_wysiwyg = "true";
defparam \rdata2_M[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N25
dffeas \rdata2_M[23] (
	.clk(CLK),
	.d(\rdata2_M~49_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_23),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[23] .is_wysiwyg = "true";
defparam \rdata2_M[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N15
dffeas \rdata2_M[24] (
	.clk(CLK),
	.d(\rdata2_M~51_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_24),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[24] .is_wysiwyg = "true";
defparam \rdata2_M[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N13
dffeas \rdata2_M[25] (
	.clk(CLK),
	.d(\rdata2_M~53_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_25),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[25] .is_wysiwyg = "true";
defparam \rdata2_M[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N7
dffeas \rdata2_M[26] (
	.clk(CLK),
	.d(\rdata2_M~55_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_26),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[26] .is_wysiwyg = "true";
defparam \rdata2_M[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N1
dffeas \rdata2_M[27] (
	.clk(CLK),
	.d(\rdata2_M~57_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_27),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[27] .is_wysiwyg = "true";
defparam \rdata2_M[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N17
dffeas \rdata2_M[28] (
	.clk(CLK),
	.d(\rdata2_M~59_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_28),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[28] .is_wysiwyg = "true";
defparam \rdata2_M[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N1
dffeas \rdata2_M[29] (
	.clk(CLK),
	.d(\rdata2_M~61_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_29),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[29] .is_wysiwyg = "true";
defparam \rdata2_M[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N23
dffeas \rdata2_M[30] (
	.clk(CLK),
	.d(\rdata2_M~63_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_30),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[30] .is_wysiwyg = "true";
defparam \rdata2_M[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N1
dffeas \rdata2_M[31] (
	.clk(CLK),
	.d(\rdata2_M~65_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\wsel_M~0_combout ),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_M_31),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_M[31] .is_wysiwyg = "true";
defparam \rdata2_M[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N25
dffeas \porto_M[1] (
	.clk(CLK),
	.d(\porto_M~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_1),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[1] .is_wysiwyg = "true";
defparam \porto_M[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N1
dffeas dWEN_M(
	.clk(CLK),
	.d(\dWEN_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dWEN_M1),
	.prn(vcc));
// synopsys translate_off
defparam dWEN_M.is_wysiwyg = "true";
defparam dWEN_M.power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N31
dffeas dREN_M(
	.clk(CLK),
	.d(\dREN_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dREN_M1),
	.prn(vcc));
// synopsys translate_off
defparam dREN_M.is_wysiwyg = "true";
defparam dREN_M.power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N1
dffeas \porto_M[0] (
	.clk(CLK),
	.d(\porto_M~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_0),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[0] .is_wysiwyg = "true";
defparam \porto_M[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N9
dffeas \porto_M[3] (
	.clk(CLK),
	.d(\porto_M~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_3),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[3] .is_wysiwyg = "true";
defparam \porto_M[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N1
dffeas \porto_M[2] (
	.clk(CLK),
	.d(\porto_M~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_2),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[2] .is_wysiwyg = "true";
defparam \porto_M[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N1
dffeas \porto_M[5] (
	.clk(CLK),
	.d(\porto_M~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_5),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[5] .is_wysiwyg = "true";
defparam \porto_M[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N1
dffeas \porto_M[4] (
	.clk(CLK),
	.d(\porto_M~36_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_4),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[4] .is_wysiwyg = "true";
defparam \porto_M[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N21
dffeas \porto_M[7] (
	.clk(CLK),
	.d(\porto_M~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_7),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[7] .is_wysiwyg = "true";
defparam \porto_M[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N9
dffeas \porto_M[6] (
	.clk(CLK),
	.d(\porto_M~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_6),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[6] .is_wysiwyg = "true";
defparam \porto_M[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N13
dffeas \porto_M[9] (
	.clk(CLK),
	.d(\porto_M~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_9),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[9] .is_wysiwyg = "true";
defparam \porto_M[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N17
dffeas \porto_M[8] (
	.clk(CLK),
	.d(\porto_M~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_8),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[8] .is_wysiwyg = "true";
defparam \porto_M[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N1
dffeas \porto_M[11] (
	.clk(CLK),
	.d(\porto_M~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_11),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[11] .is_wysiwyg = "true";
defparam \porto_M[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N21
dffeas \porto_M[10] (
	.clk(CLK),
	.d(\porto_M~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_10),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[10] .is_wysiwyg = "true";
defparam \porto_M[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N19
dffeas \porto_M[13] (
	.clk(CLK),
	.d(\porto_M~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_13),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[13] .is_wysiwyg = "true";
defparam \porto_M[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N23
dffeas \porto_M[12] (
	.clk(CLK),
	.d(\porto_M~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_12),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[12] .is_wysiwyg = "true";
defparam \porto_M[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N19
dffeas \porto_M[15] (
	.clk(CLK),
	.d(\porto_M~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_15),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[15] .is_wysiwyg = "true";
defparam \porto_M[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N29
dffeas \porto_M[14] (
	.clk(CLK),
	.d(\porto_M~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_14),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[14] .is_wysiwyg = "true";
defparam \porto_M[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N11
dffeas \porto_M[17] (
	.clk(CLK),
	.d(\porto_M~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_17),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[17] .is_wysiwyg = "true";
defparam \porto_M[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N21
dffeas \porto_M[16] (
	.clk(CLK),
	.d(\porto_M~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_16),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[16] .is_wysiwyg = "true";
defparam \porto_M[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y28_N17
dffeas \porto_M[19] (
	.clk(CLK),
	.d(\porto_M~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_19),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[19] .is_wysiwyg = "true";
defparam \porto_M[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N19
dffeas \porto_M[18] (
	.clk(CLK),
	.d(\porto_M~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_18),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[18] .is_wysiwyg = "true";
defparam \porto_M[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y28_N7
dffeas \porto_M[21] (
	.clk(CLK),
	.d(\porto_M~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_21),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[21] .is_wysiwyg = "true";
defparam \porto_M[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N15
dffeas \porto_M[20] (
	.clk(CLK),
	.d(\porto_M~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_20),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[20] .is_wysiwyg = "true";
defparam \porto_M[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N29
dffeas \porto_M[23] (
	.clk(CLK),
	.d(\porto_M~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_23),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[23] .is_wysiwyg = "true";
defparam \porto_M[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N15
dffeas \porto_M[22] (
	.clk(CLK),
	.d(\porto_M~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_22),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[22] .is_wysiwyg = "true";
defparam \porto_M[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N21
dffeas \porto_M[25] (
	.clk(CLK),
	.d(\porto_M~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_25),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[25] .is_wysiwyg = "true";
defparam \porto_M[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N17
dffeas \porto_M[24] (
	.clk(CLK),
	.d(\porto_M~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_24),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[24] .is_wysiwyg = "true";
defparam \porto_M[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N19
dffeas \porto_M[27] (
	.clk(CLK),
	.d(\porto_M~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_27),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[27] .is_wysiwyg = "true";
defparam \porto_M[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N31
dffeas \porto_M[26] (
	.clk(CLK),
	.d(\porto_M~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_26),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[26] .is_wysiwyg = "true";
defparam \porto_M[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N17
dffeas \porto_M[29] (
	.clk(CLK),
	.d(\porto_M~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_29),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[29] .is_wysiwyg = "true";
defparam \porto_M[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N15
dffeas \porto_M[28] (
	.clk(CLK),
	.d(\porto_M~32_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_28),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[28] .is_wysiwyg = "true";
defparam \porto_M[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N31
dffeas \porto_M[31] (
	.clk(CLK),
	.d(\porto_M~33_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_31),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[31] .is_wysiwyg = "true";
defparam \porto_M[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N3
dffeas \porto_M[30] (
	.clk(CLK),
	.d(\porto_M~34_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_M_30),
	.prn(vcc));
// synopsys translate_off
defparam \porto_M[30] .is_wysiwyg = "true";
defparam \porto_M[30] .power_up = "low";
// synopsys translate_on

// Location: DDIOOUTCELL_X60_Y0_N11
dffeas halt_WB(
	.clk(CLK),
	.d(\halt_M~q ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(halt_WB1),
	.prn(vcc));
// synopsys translate_off
defparam halt_WB.is_wysiwyg = "true";
defparam halt_WB.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N26
cycloneive_lcell_comb \instruction_D~68 (
// Equation(s):
// \instruction_D~68_combout  = (iwait & (\branch_or_jump~1_combout  & ramiframload_27))

	.dataa(iwait),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\dpif.dmemload [27]),
	.cin(gnd),
	.combout(\instruction_D~68_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~68 .lut_mask = 16'hA000;
defparam \instruction_D~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N26
cycloneive_lcell_comb \ALUSrc_EX~0 (
// Equation(s):
// \ALUSrc_EX~0_combout  = ((always1 & ((!dhit) # (!fuifbubble_lw_f)))) # (!\branch_or_jump~1_combout )

	.dataa(\FORWARDING_UNIT|fuif.bubble_lw_f~2_combout ),
	.datab(dhit),
	.datac(\branch_or_jump~1_combout ),
	.datad(always1),
	.cin(gnd),
	.combout(\ALUSrc_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSrc_EX~0 .lut_mask = 16'h7F0F;
defparam \ALUSrc_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N27
dffeas \instruction_D[27] (
	.clk(CLK),
	.d(\instruction_D~68_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[27]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[27] .is_wysiwyg = "true";
defparam \instruction_D[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N10
cycloneive_lcell_comb \instruction_D~69 (
// Equation(s):
// \instruction_D~69_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_26))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(\dpif.dmemload [26]),
	.cin(gnd),
	.combout(\instruction_D~69_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~69 .lut_mask = 16'hC000;
defparam \instruction_D~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N11
dffeas \instruction_D[26] (
	.clk(CLK),
	.d(\instruction_D~69_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[26]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[26] .is_wysiwyg = "true";
defparam \instruction_D[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N20
cycloneive_lcell_comb \instruction_D~66 (
// Equation(s):
// \instruction_D~66_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_30))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(\dpif.dmemload [30]),
	.cin(gnd),
	.combout(\instruction_D~66_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~66 .lut_mask = 16'hC000;
defparam \instruction_D~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N21
dffeas \instruction_D[30] (
	.clk(CLK),
	.d(\instruction_D~66_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[30]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[30] .is_wysiwyg = "true";
defparam \instruction_D[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N28
cycloneive_lcell_comb \instruction_D~67 (
// Equation(s):
// \instruction_D~67_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_29))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(iwait),
	.datad(\dpif.dmemload [29]),
	.cin(gnd),
	.combout(\instruction_D~67_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~67 .lut_mask = 16'hA000;
defparam \instruction_D~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N29
dffeas \instruction_D[29] (
	.clk(CLK),
	.d(\instruction_D~67_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[29]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[29] .is_wysiwyg = "true";
defparam \instruction_D[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N6
cycloneive_lcell_comb \j_EX~3 (
// Equation(s):
// \j_EX~3_combout  = (!instruction_D[31] & (!instruction_D[30] & (!instruction_D[29] & \branch_or_jump~1_combout )))

	.dataa(instruction_D[31]),
	.datab(instruction_D[30]),
	.datac(instruction_D[29]),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\j_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \j_EX~3 .lut_mask = 16'h0100;
defparam \j_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N6
cycloneive_lcell_comb \j_EX~2 (
// Equation(s):
// \j_EX~2_combout  = (!instruction_D[28] & (instruction_D[27] & (!instruction_D[26] & \j_EX~3_combout )))

	.dataa(instruction_D[28]),
	.datab(instruction_D[27]),
	.datac(instruction_D[26]),
	.datad(\j_EX~3_combout ),
	.cin(gnd),
	.combout(\j_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \j_EX~2 .lut_mask = 16'h0400;
defparam \j_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N7
dffeas j_EX(
	.clk(CLK),
	.d(\j_EX~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\j_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam j_EX.is_wysiwyg = "true";
defparam j_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N10
cycloneive_lcell_comb \predicted_M~3 (
// Equation(s):
// \predicted_M~3_combout  = (always1 & (((!dREN_M1 & !dWEN_M1)) # (!fuifbubble_lw_f)))

	.dataa(dREN_M1),
	.datab(dWEN_M1),
	.datac(always1),
	.datad(\FORWARDING_UNIT|fuif.bubble_lw_f~2_combout ),
	.cin(gnd),
	.combout(\predicted_M~3_combout ),
	.cout());
// synopsys translate_off
defparam \predicted_M~3 .lut_mask = 16'h10F0;
defparam \predicted_M~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N12
cycloneive_lcell_comb \j_M~0 (
// Equation(s):
// \j_M~0_combout  = (\branch_or_jump~1_combout  & (\j_EX~q  & \predicted_M~3_combout ))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(\j_EX~q ),
	.datad(\predicted_M~3_combout ),
	.cin(gnd),
	.combout(\j_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \j_M~0 .lut_mask = 16'hA000;
defparam \j_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N13
dffeas j_M(
	.clk(CLK),
	.d(\j_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\j_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam j_M.is_wysiwyg = "true";
defparam j_M.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N8
cycloneive_lcell_comb \en_EX~0 (
// Equation(s):
// \en_EX~0_combout  = (\nRST~input_o  & ((!always0) # (!LessThan1)))

	.dataa(gnd),
	.datab(LessThan1),
	.datac(nRST),
	.datad(always0),
	.cin(gnd),
	.combout(\en_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \en_EX~0 .lut_mask = 16'h30F0;
defparam \en_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N14
cycloneive_lcell_comb \wsel_M~0 (
// Equation(s):
// \wsel_M~0_combout  = ((fuifbubble_lw_f & (dhit & always1))) # (!\branch_or_jump~1_combout )

	.dataa(\FORWARDING_UNIT|fuif.bubble_lw_f~2_combout ),
	.datab(dhit),
	.datac(\branch_or_jump~1_combout ),
	.datad(always1),
	.cin(gnd),
	.combout(\wsel_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \wsel_M~0 .lut_mask = 16'h8F0F;
defparam \wsel_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N14
cycloneive_lcell_comb \jal_M~0 (
// Equation(s):
// \jal_M~0_combout  = (\jal_EX~q  & (!\en_EX~0_combout  & !\wsel_M~0_combout ))

	.dataa(\jal_EX~q ),
	.datab(gnd),
	.datac(\en_EX~0_combout ),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\jal_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \jal_M~0 .lut_mask = 16'h000A;
defparam \jal_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N15
dffeas jal_M(
	.clk(CLK),
	.d(\jal_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\jal_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam jal_M.is_wysiwyg = "true";
defparam jal_M.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N2
cycloneive_lcell_comb \branch_or_jump~0 (
// Equation(s):
// \branch_or_jump~0_combout  = (!\j_M~q  & !\jal_M~q )

	.dataa(gnd),
	.datab(gnd),
	.datac(\j_M~q ),
	.datad(\jal_M~q ),
	.cin(gnd),
	.combout(\branch_or_jump~0_combout ),
	.cout());
// synopsys translate_off
defparam \branch_or_jump~0 .lut_mask = 16'h000F;
defparam \branch_or_jump~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N0
cycloneive_lcell_comb \predicted_M~2 (
// Equation(s):
// \predicted_M~2_combout  = (\predicted_EX~q  & ((\predicted_M~3_combout ) # ((\en_EX~0_combout  & \predicted_M~q )))) # (!\predicted_EX~q  & (\en_EX~0_combout  & (\predicted_M~q )))

	.dataa(\predicted_EX~q ),
	.datab(\en_EX~0_combout ),
	.datac(\predicted_M~q ),
	.datad(\predicted_M~3_combout ),
	.cin(gnd),
	.combout(\predicted_M~2_combout ),
	.cout());
// synopsys translate_off
defparam \predicted_M~2 .lut_mask = 16'hEAC0;
defparam \predicted_M~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N1
dffeas predicted_M(
	.clk(CLK),
	.d(\predicted_M~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\predicted_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam predicted_M.is_wysiwyg = "true";
defparam predicted_M.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N20
cycloneive_lcell_comb \beq_M~0 (
// Equation(s):
// \beq_M~0_combout  = (\beq_EX~q  & !\wsel_M~0_combout )

	.dataa(\beq_EX~q ),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\beq_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \beq_M~0 .lut_mask = 16'h0A0A;
defparam \beq_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N30
cycloneive_lcell_comb \always4~3 (
// Equation(s):
// \always4~3_combout  = (((LessThan1 & always0)) # (!\nRST~input_o )) # (!\branch_or_jump~1_combout )

	.dataa(LessThan1),
	.datab(\branch_or_jump~1_combout ),
	.datac(nRST),
	.datad(always0),
	.cin(gnd),
	.combout(\always4~3_combout ),
	.cout());
// synopsys translate_off
defparam \always4~3 .lut_mask = 16'hBF3F;
defparam \always4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N21
dffeas beq_M(
	.clk(CLK),
	.d(\beq_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\beq_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam beq_M.is_wysiwyg = "true";
defparam beq_M.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N8
cycloneive_lcell_comb \zero_M~7 (
// Equation(s):
// \zero_M~7_combout  = (!Selector17 & (!Selector13 & (!Selector14 & !Selector18)))

	.dataa(\ALU|Selector17~8_combout ),
	.datab(\ALU|Selector13~8_combout ),
	.datac(\ALU|Selector14~7_combout ),
	.datad(\ALU|Selector18~7_combout ),
	.cin(gnd),
	.combout(\zero_M~7_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~7 .lut_mask = 16'h0001;
defparam \zero_M~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N30
cycloneive_lcell_comb \zero_M~8 (
// Equation(s):
// \zero_M~8_combout  = (!Selector23 & (!Selector11 & (\zero_M~7_combout  & !Selector121)))

	.dataa(\ALU|Selector23~8_combout ),
	.datab(\ALU|Selector11~8_combout ),
	.datac(\zero_M~7_combout ),
	.datad(\ALU|Selector12~18_combout ),
	.cin(gnd),
	.combout(\zero_M~8_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~8 .lut_mask = 16'h0010;
defparam \zero_M~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N22
cycloneive_lcell_comb \zero_M~9 (
// Equation(s):
// \zero_M~9_combout  = (Selector21) # ((Selector19) # ((ShiftLeft0 & Selector16)))

	.dataa(\ALU|ShiftLeft0~57_combout ),
	.datab(\ALU|Selector16~3_combout ),
	.datac(\ALU|Selector21~7_combout ),
	.datad(\ALU|Selector19~6_combout ),
	.cin(gnd),
	.combout(\zero_M~9_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~9 .lut_mask = 16'hFFF8;
defparam \zero_M~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N12
cycloneive_lcell_comb \zero_M~10 (
// Equation(s):
// \zero_M~10_combout  = (Selector10) # ((\zero_M~9_combout ) # ((Selector9) # (Selector20)))

	.dataa(\ALU|Selector10~8_combout ),
	.datab(\zero_M~9_combout ),
	.datac(\ALU|Selector9~8_combout ),
	.datad(\ALU|Selector20~8_combout ),
	.cin(gnd),
	.combout(\zero_M~10_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~10 .lut_mask = 16'hFFFE;
defparam \zero_M~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N14
cycloneive_lcell_comb \zero_M~11 (
// Equation(s):
// \zero_M~11_combout  = (!Selector22 & (!Selector1 & (\zero_M~8_combout  & !\zero_M~10_combout )))

	.dataa(\ALU|Selector22~8_combout ),
	.datab(\ALU|Selector1~9_combout ),
	.datac(\zero_M~8_combout ),
	.datad(\zero_M~10_combout ),
	.cin(gnd),
	.combout(\zero_M~11_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~11 .lut_mask = 16'h0010;
defparam \zero_M~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N6
cycloneive_lcell_comb \zero_M~0 (
// Equation(s):
// \zero_M~0_combout  = (!Selector61 & (!Selector64 & (!Selector6 & !Selector24)))

	.dataa(\ALU|Selector6~5_combout ),
	.datab(\ALU|Selector6~9_combout ),
	.datac(\ALU|Selector6~0_combout ),
	.datad(\ALU|Selector24~8_combout ),
	.cin(gnd),
	.combout(\zero_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~0 .lut_mask = 16'h0001;
defparam \zero_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N26
cycloneive_lcell_comb \zero_M~1 (
// Equation(s):
// \zero_M~1_combout  = (!Selector25 & (!Selector26 & (!Selector273 & \zero_M~0_combout )))

	.dataa(\ALU|Selector25~7_combout ),
	.datab(\ALU|Selector26~6_combout ),
	.datac(\ALU|Selector27~7_combout ),
	.datad(\zero_M~0_combout ),
	.cin(gnd),
	.combout(\zero_M~1_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~1 .lut_mask = 16'h0100;
defparam \zero_M~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N4
cycloneive_lcell_comb \zero_M~2 (
// Equation(s):
// \zero_M~2_combout  = (!Selector7 & (!Selector63 & (\zero_M~1_combout  & !Selector15)))

	.dataa(\ALU|Selector7~7_combout ),
	.datab(\ALU|Selector6~8_combout ),
	.datac(\zero_M~1_combout ),
	.datad(\ALU|Selector15~11_combout ),
	.cin(gnd),
	.combout(\zero_M~2_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~2 .lut_mask = 16'h0010;
defparam \zero_M~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N22
cycloneive_lcell_comb \zero_M~3 (
// Equation(s):
// \zero_M~3_combout  = (!\wsel_M~0_combout  & (!Selector4 & (!Selector29 & !Selector5)))

	.dataa(\wsel_M~0_combout ),
	.datab(\ALU|Selector4~12_combout ),
	.datac(\ALU|Selector29~10_combout ),
	.datad(\ALU|Selector5~7_combout ),
	.cin(gnd),
	.combout(\zero_M~3_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~3 .lut_mask = 16'h0001;
defparam \zero_M~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N28
cycloneive_lcell_comb \zero_M~4 (
// Equation(s):
// \zero_M~4_combout  = (!Selector28 & (!Selector3 & (\zero_M~3_combout  & !Selector2)))

	.dataa(\ALU|Selector28~10_combout ),
	.datab(\ALU|Selector3~9_combout ),
	.datac(\zero_M~3_combout ),
	.datad(\ALU|Selector2~11_combout ),
	.cin(gnd),
	.combout(\zero_M~4_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~4 .lut_mask = 16'h0010;
defparam \zero_M~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N2
cycloneive_lcell_comb \zero_M~6 (
// Equation(s):
// \zero_M~6_combout  = (!\zero_M~5_combout  & (!Selector8 & (\zero_M~2_combout  & \zero_M~4_combout )))

	.dataa(\zero_M~5_combout ),
	.datab(\ALU|Selector8~7_combout ),
	.datac(\zero_M~2_combout ),
	.datad(\zero_M~4_combout ),
	.cin(gnd),
	.combout(\zero_M~6_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~6 .lut_mask = 16'h1000;
defparam \zero_M~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N24
cycloneive_lcell_comb \zero_M~12 (
// Equation(s):
// \zero_M~12_combout  = (!Selector01 & (!Selector313 & (\zero_M~11_combout  & \zero_M~6_combout )))

	.dataa(\ALU|Selector0~27_combout ),
	.datab(\ALU|Selector31~9_combout ),
	.datac(\zero_M~11_combout ),
	.datad(\zero_M~6_combout ),
	.cin(gnd),
	.combout(\zero_M~12_combout ),
	.cout());
// synopsys translate_off
defparam \zero_M~12 .lut_mask = 16'h1000;
defparam \zero_M~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N25
dffeas zero_M(
	.clk(CLK),
	.d(\zero_M~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\zero_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam zero_M.is_wysiwyg = "true";
defparam zero_M.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N16
cycloneive_lcell_comb \branch_taken~0 (
// Equation(s):
// \branch_taken~0_combout  = (\zero_M~q  & ((\beq_M~q ))) # (!\zero_M~q  & (\bne_M~q ))

	.dataa(\bne_M~q ),
	.datab(\beq_M~q ),
	.datac(gnd),
	.datad(\zero_M~q ),
	.cin(gnd),
	.combout(\branch_taken~0_combout ),
	.cout());
// synopsys translate_off
defparam \branch_taken~0 .lut_mask = 16'hCCAA;
defparam \branch_taken~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N4
cycloneive_lcell_comb \branch_or_jump~1 (
// Equation(s):
// \branch_or_jump~1_combout  = (!\jr_M~q  & (\branch_or_jump~0_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\jr_M~q ),
	.datab(\branch_or_jump~0_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\branch_or_jump~1_combout ),
	.cout());
// synopsys translate_off
defparam \branch_or_jump~1 .lut_mask = 16'h4004;
defparam \branch_or_jump~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N0
cycloneive_lcell_comb \pc_plus_4_D~1 (
// Equation(s):
// \pc_plus_4_D~1_combout  = (pc_out_0 & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(iwait),
	.datab(gnd),
	.datac(pc_out_0),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~1_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~1 .lut_mask = 16'hA0F0;
defparam \pc_plus_4_D~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N1
dffeas \pc_plus_4_D[0] (
	.clk(CLK),
	.d(\pc_plus_4_D~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[0]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[0] .is_wysiwyg = "true";
defparam \pc_plus_4_D[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N22
cycloneive_lcell_comb \branch_or_jump~2 (
// Equation(s):
// \branch_or_jump~2_combout  = (!\jr_M~q  & (!\j_M~q  & !\jal_M~q ))

	.dataa(\jr_M~q ),
	.datab(gnd),
	.datac(\j_M~q ),
	.datad(\jal_M~q ),
	.cin(gnd),
	.combout(\branch_or_jump~2_combout ),
	.cout());
// synopsys translate_off
defparam \branch_or_jump~2 .lut_mask = 16'h0005;
defparam \branch_or_jump~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N16
cycloneive_lcell_comb \pc_plus_4_EX~1 (
// Equation(s):
// \pc_plus_4_EX~1_combout  = (pc_plus_4_D[0] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(pc_plus_4_D[0]),
	.datac(\branch_taken~0_combout ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~1 .lut_mask = 16'h8400;
defparam \pc_plus_4_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N17
dffeas \pc_plus_4_EX[0] (
	.clk(CLK),
	.d(\pc_plus_4_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[0]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[0] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N16
cycloneive_lcell_comb \pc_plus_4_M~1 (
// Equation(s):
// \pc_plus_4_M~1_combout  = (pc_plus_4_EX[0] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[0]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~1_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~1 .lut_mask = 16'h00CC;
defparam \pc_plus_4_M~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N17
dffeas \pc_plus_4_M[0] (
	.clk(CLK),
	.d(\pc_plus_4_M~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[0]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[0] .is_wysiwyg = "true";
defparam \pc_plus_4_M[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N4
cycloneive_lcell_comb \pc_plus_4_WB[0]~feeder (
// Equation(s):
// \pc_plus_4_WB[0]~feeder_combout  = pc_plus_4_M[0]

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pc_plus_4_M[0]),
	.cin(gnd),
	.combout(\pc_plus_4_WB[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_WB[0]~feeder .lut_mask = 16'hFF00;
defparam \pc_plus_4_WB[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N8
cycloneive_lcell_comb \halt_M~0 (
// Equation(s):
// \halt_M~0_combout  = (\cu_halt_EX~q  & !\wsel_M~0_combout )

	.dataa(\cu_halt_EX~q ),
	.datab(\wsel_M~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\halt_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \halt_M~0 .lut_mask = 16'h2222;
defparam \halt_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N9
dffeas halt_M(
	.clk(CLK),
	.d(\halt_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\halt_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam halt_M.is_wysiwyg = "true";
defparam halt_M.power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N9
dffeas \halt_WB~_Duplicate_1 (
	.clk(CLK),
	.d(gnd),
	.asdata(\halt_M~q ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\halt_WB~_Duplicate_1_q ),
	.prn(vcc));
// synopsys translate_off
defparam \halt_WB~_Duplicate_1 .is_wysiwyg = "true";
defparam \halt_WB~_Duplicate_1 .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N8
cycloneive_lcell_comb \always4~2 (
// Equation(s):
// \always4~2_combout  = (!\halt_WB~_Duplicate_1_q  & ((!\en_EX~0_combout ) # (!\branch_or_jump~1_combout )))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(\halt_WB~_Duplicate_1_q ),
	.datad(\en_EX~0_combout ),
	.cin(gnd),
	.combout(\always4~2_combout ),
	.cout());
// synopsys translate_off
defparam \always4~2 .lut_mask = 16'h050F;
defparam \always4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N5
dffeas \pc_plus_4_WB[0] (
	.clk(CLK),
	.d(\pc_plus_4_WB[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[0]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[0] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N14
cycloneive_lcell_comb \lui_M~0 (
// Equation(s):
// \lui_M~0_combout  = (\lui_EX~q  & !\wsel_M~0_combout )

	.dataa(\lui_EX~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\lui_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \lui_M~0 .lut_mask = 16'h00AA;
defparam \lui_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N15
dffeas lui_M(
	.clk(CLK),
	.d(\lui_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\lui_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam lui_M.is_wysiwyg = "true";
defparam lui_M.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N29
dffeas lui_WB(
	.clk(CLK),
	.d(gnd),
	.asdata(\lui_M~q ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\lui_WB~q ),
	.prn(vcc));
// synopsys translate_off
defparam lui_WB.is_wysiwyg = "true";
defparam lui_WB.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N17
dffeas \dmemload_WB[0] (
	.clk(CLK),
	.d(\dpif.dmemload [0]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[0]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[0] .is_wysiwyg = "true";
defparam \dmemload_WB[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N25
dffeas \porto_WB[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_0),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[0]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[0] .is_wysiwyg = "true";
defparam \porto_WB[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N6
cycloneive_lcell_comb \jal_WB~feeder (
// Equation(s):
// \jal_WB~feeder_combout  = \jal_M~q 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\jal_M~q ),
	.cin(gnd),
	.combout(\jal_WB~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \jal_WB~feeder .lut_mask = 16'hFF00;
defparam \jal_WB~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N7
dffeas jal_WB(
	.clk(CLK),
	.d(\jal_WB~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\jal_WB~q ),
	.prn(vcc));
// synopsys translate_off
defparam jal_WB.is_wysiwyg = "true";
defparam jal_WB.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N24
cycloneive_lcell_comb \wdat_WB[0]~60 (
// Equation(s):
// \wdat_WB[0]~60_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[0])) # (!\memToReg_WB~q  & ((porto_WB[0])))))

	.dataa(\memToReg_WB~q ),
	.datab(dmemload_WB[0]),
	.datac(porto_WB[0]),
	.datad(\jal_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[0]~60_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[0]~60 .lut_mask = 16'h00D8;
defparam \wdat_WB[0]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N26
cycloneive_lcell_comb \wdat_WB[0]~61 (
// Equation(s):
// \wdat_WB[0]~61_combout  = (!\lui_WB~q  & ((\wdat_WB[0]~60_combout ) # ((\jal_WB~q  & pc_plus_4_WB[0]))))

	.dataa(\jal_WB~q ),
	.datab(pc_plus_4_WB[0]),
	.datac(\lui_WB~q ),
	.datad(\wdat_WB[0]~60_combout ),
	.cin(gnd),
	.combout(\wdat_WB[0]~61_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[0]~61 .lut_mask = 16'h0F08;
defparam \wdat_WB[0]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N12
cycloneive_lcell_comb \instruction_D~65 (
// Equation(s):
// \instruction_D~65_combout  = (\branch_or_jump~1_combout  & (ramiframload_28 & iwait))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(\dpif.dmemload [28]),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~65_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~65 .lut_mask = 16'hC000;
defparam \instruction_D~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N13
dffeas \instruction_D[28] (
	.clk(CLK),
	.d(\instruction_D~65_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[28]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[28] .is_wysiwyg = "true";
defparam \instruction_D[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N2
cycloneive_lcell_comb \instruction_D~64 (
// Equation(s):
// \instruction_D~64_combout  = (\branch_or_jump~1_combout  & (ramiframload_31 & iwait))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(\dpif.dmemload [31]),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~64_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~64 .lut_mask = 16'hC000;
defparam \instruction_D~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N3
dffeas \instruction_D[31] (
	.clk(CLK),
	.d(\instruction_D~64_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[31]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[31] .is_wysiwyg = "true";
defparam \instruction_D[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N26
cycloneive_lcell_comb \dWEN_EX~0 (
// Equation(s):
// \dWEN_EX~0_combout  = (\lui_EX~0_combout  & (instruction_D[29] & (!instruction_D[28] & instruction_D[31])))

	.dataa(\lui_EX~0_combout ),
	.datab(instruction_D[29]),
	.datac(instruction_D[28]),
	.datad(instruction_D[31]),
	.cin(gnd),
	.combout(\dWEN_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \dWEN_EX~0 .lut_mask = 16'h0800;
defparam \dWEN_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N27
dffeas dWEN_EX(
	.clk(CLK),
	.d(\dWEN_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\dWEN_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam dWEN_EX.is_wysiwyg = "true";
defparam dWEN_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N26
cycloneive_lcell_comb \rdata2_M[16]~0 (
// Equation(s):
// \rdata2_M[16]~0_combout  = (\dWEN_EX~q  & ((Equal0 & (dREN_M1)) # (!Equal0 & ((fuifforward_B_1)))))

	.dataa(\FORWARDING_UNIT|Equal0~2_combout ),
	.datab(\dWEN_EX~q ),
	.datac(dREN_M1),
	.datad(\FORWARDING_UNIT|fuif.forward_B[1]~3_combout ),
	.cin(gnd),
	.combout(\rdata2_M[16]~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M[16]~0 .lut_mask = 16'hC480;
defparam \rdata2_M[16]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N12
cycloneive_lcell_comb \rdata2_M[16]~1 (
// Equation(s):
// \rdata2_M[16]~1_combout  = (\dWEN_EX~q  & ((Equal0 & (!dREN_M1)) # (!Equal0 & ((fuifforward_B_1)))))

	.dataa(\FORWARDING_UNIT|Equal0~2_combout ),
	.datab(\dWEN_EX~q ),
	.datac(dREN_M1),
	.datad(\FORWARDING_UNIT|fuif.forward_B[1]~3_combout ),
	.cin(gnd),
	.combout(\rdata2_M[16]~1_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M[16]~1 .lut_mask = 16'h4C08;
defparam \rdata2_M[16]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N12
cycloneive_lcell_comb \sw_forwarding_output~27 (
// Equation(s):
// \sw_forwarding_output~27_combout  = (porto_M_0 & !\lui_M~q )

	.dataa(gnd),
	.datab(porto_M_0),
	.datac(\lui_M~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sw_forwarding_output~27_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~27 .lut_mask = 16'h0C0C;
defparam \sw_forwarding_output~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N14
cycloneive_lcell_comb \rdata2_M~2 (
// Equation(s):
// \rdata2_M~2_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & ((\rdata2_M[16]~1_combout  & ((\sw_forwarding_output~27_combout ))) # (!\rdata2_M[16]~1_combout  & (rdata2_EX[0]))))

	.dataa(rdata2_EX[0]),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\sw_forwarding_output~27_combout ),
	.cin(gnd),
	.combout(\rdata2_M~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~2 .lut_mask = 16'hF2C2;
defparam \rdata2_M~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N4
cycloneive_lcell_comb \rdata2_M~3 (
// Equation(s):
// \rdata2_M~3_combout  = (\rdata2_M[16]~0_combout  & ((\rdata2_M~2_combout  & (\wdat_WB[0]~61_combout )) # (!\rdata2_M~2_combout  & ((ramiframload_0))))) # (!\rdata2_M[16]~0_combout  & (((\rdata2_M~2_combout ))))

	.dataa(\wdat_WB[0]~61_combout ),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\rdata2_M~2_combout ),
	.datad(\dpif.dmemload [0]),
	.cin(gnd),
	.combout(\rdata2_M~3_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~3 .lut_mask = 16'hBCB0;
defparam \rdata2_M~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N2
cycloneive_lcell_comb \sw_forwarding_output~28 (
// Equation(s):
// \sw_forwarding_output~28_combout  = (porto_M_1 & !\lui_M~q )

	.dataa(gnd),
	.datab(gnd),
	.datac(porto_M_1),
	.datad(\lui_M~q ),
	.cin(gnd),
	.combout(\sw_forwarding_output~28_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~28 .lut_mask = 16'h00F0;
defparam \sw_forwarding_output~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N15
dffeas \dmemload_WB[1] (
	.clk(CLK),
	.d(\dpif.dmemload [1]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[1]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[1] .is_wysiwyg = "true";
defparam \dmemload_WB[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N3
dffeas \porto_WB[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_1),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[1]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[1] .is_wysiwyg = "true";
defparam \porto_WB[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N14
cycloneive_lcell_comb \lui_EX~0 (
// Equation(s):
// \lui_EX~0_combout  = (instruction_D[26] & (\branch_or_jump~1_combout  & (!instruction_D[30] & instruction_D[27])))

	.dataa(instruction_D[26]),
	.datab(\branch_or_jump~1_combout ),
	.datac(instruction_D[30]),
	.datad(instruction_D[27]),
	.cin(gnd),
	.combout(\lui_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \lui_EX~0 .lut_mask = 16'h0800;
defparam \lui_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N14
cycloneive_lcell_comb \MemToReg_EX~2 (
// Equation(s):
// \MemToReg_EX~2_combout  = (instruction_D[31] & (!instruction_D[29] & (\lui_EX~0_combout  & !instruction_D[28])))

	.dataa(instruction_D[31]),
	.datab(instruction_D[29]),
	.datac(\lui_EX~0_combout ),
	.datad(instruction_D[28]),
	.cin(gnd),
	.combout(\MemToReg_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \MemToReg_EX~2 .lut_mask = 16'h0020;
defparam \MemToReg_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N15
dffeas MemToReg_EX(
	.clk(CLK),
	.d(\MemToReg_EX~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\MemToReg_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam MemToReg_EX.is_wysiwyg = "true";
defparam MemToReg_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N22
cycloneive_lcell_comb \memToReg_M~0 (
// Equation(s):
// \memToReg_M~0_combout  = (!\wsel_M~0_combout  & \MemToReg_EX~q )

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(\MemToReg_EX~q ),
	.cin(gnd),
	.combout(\memToReg_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \memToReg_M~0 .lut_mask = 16'h0F00;
defparam \memToReg_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N23
dffeas memToReg_M(
	.clk(CLK),
	.d(\memToReg_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\memToReg_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam memToReg_M.is_wysiwyg = "true";
defparam memToReg_M.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N31
dffeas memToReg_WB(
	.clk(CLK),
	.d(gnd),
	.asdata(\memToReg_M~q ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\memToReg_WB~q ),
	.prn(vcc));
// synopsys translate_off
defparam memToReg_WB.is_wysiwyg = "true";
defparam memToReg_WB.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N2
cycloneive_lcell_comb \wdat_WB[1]~58 (
// Equation(s):
// \wdat_WB[1]~58_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[1])) # (!\memToReg_WB~q  & ((porto_WB[1])))))

	.dataa(\jal_WB~q ),
	.datab(dmemload_WB[1]),
	.datac(porto_WB[1]),
	.datad(\memToReg_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[1]~58_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[1]~58 .lut_mask = 16'h4450;
defparam \wdat_WB[1]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N6
cycloneive_lcell_comb \pc_plus_4_M~0 (
// Equation(s):
// \pc_plus_4_M~0_combout  = (pc_plus_4_EX[1] & !\wsel_M~0_combout )

	.dataa(pc_plus_4_EX[1]),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_plus_4_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~0 .lut_mask = 16'h0A0A;
defparam \pc_plus_4_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N7
dffeas \pc_plus_4_M[1] (
	.clk(CLK),
	.d(\pc_plus_4_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[1]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[1] .is_wysiwyg = "true";
defparam \pc_plus_4_M[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N11
dffeas \pc_plus_4_WB[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[1]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[1]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[1] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N16
cycloneive_lcell_comb \wdat_WB[1]~59 (
// Equation(s):
// \wdat_WB[1]~59_combout  = (!\lui_WB~q  & ((\wdat_WB[1]~58_combout ) # ((\jal_WB~q  & pc_plus_4_WB[1]))))

	.dataa(\lui_WB~q ),
	.datab(\jal_WB~q ),
	.datac(\wdat_WB[1]~58_combout ),
	.datad(pc_plus_4_WB[1]),
	.cin(gnd),
	.combout(\wdat_WB[1]~59_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[1]~59 .lut_mask = 16'h5450;
defparam \wdat_WB[1]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N28
cycloneive_lcell_comb \rdata2_M~4 (
// Equation(s):
// \rdata2_M~4_combout  = (\rdata2_M[16]~0_combout  & (((ramiframload_1) # (\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[1] & ((!\rdata2_M[16]~1_combout ))))

	.dataa(rdata2_EX[1]),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\dpif.dmemload [1]),
	.datad(\rdata2_M[16]~1_combout ),
	.cin(gnd),
	.combout(\rdata2_M~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~4 .lut_mask = 16'hCCE2;
defparam \rdata2_M~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N8
cycloneive_lcell_comb \rdata2_M~5 (
// Equation(s):
// \rdata2_M~5_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~4_combout  & ((\wdat_WB[1]~59_combout ))) # (!\rdata2_M~4_combout  & (\sw_forwarding_output~28_combout )))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~4_combout ))))

	.dataa(\rdata2_M[16]~1_combout ),
	.datab(\sw_forwarding_output~28_combout ),
	.datac(\wdat_WB[1]~59_combout ),
	.datad(\rdata2_M~4_combout ),
	.cin(gnd),
	.combout(\rdata2_M~5_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~5 .lut_mask = 16'hF588;
defparam \rdata2_M~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N2
cycloneive_lcell_comb \pc_plus_4[2]~0 (
// Equation(s):
// \pc_plus_4[2]~0_combout  = pc_out_2 $ (VCC)
// \pc_plus_4[2]~1  = CARRY(pc_out_2)

	.dataa(gnd),
	.datab(pc_out_2),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\pc_plus_4[2]~0_combout ),
	.cout(\pc_plus_4[2]~1 ));
// synopsys translate_off
defparam \pc_plus_4[2]~0 .lut_mask = 16'h33CC;
defparam \pc_plus_4[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N28
cycloneive_lcell_comb \pc_plus_4_D~3 (
// Equation(s):
// \pc_plus_4_D~3_combout  = (\pc_plus_4[2]~0_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\branch_or_jump~1_combout ),
	.datab(\pc_plus_4[2]~0_combout ),
	.datac(gnd),
	.datad(iwait),
	.cin(gnd),
	.combout(\pc_plus_4_D~3_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~3 .lut_mask = 16'hCC44;
defparam \pc_plus_4_D~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N29
dffeas \pc_plus_4_D[2] (
	.clk(CLK),
	.d(\pc_plus_4_D~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[2]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[2] .is_wysiwyg = "true";
defparam \pc_plus_4_D[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N30
cycloneive_lcell_comb \pc_plus_4_EX~3 (
// Equation(s):
// \pc_plus_4_EX~3_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[2] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_D[2]),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~3 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N31
dffeas \pc_plus_4_EX[2] (
	.clk(CLK),
	.d(\pc_plus_4_EX~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[2]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[2] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N12
cycloneive_lcell_comb \pc_plus_4_M~3 (
// Equation(s):
// \pc_plus_4_M~3_combout  = (pc_plus_4_EX[2] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_plus_4_EX[2]),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~3_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~3 .lut_mask = 16'h00F0;
defparam \pc_plus_4_M~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y39_N13
dffeas \pc_plus_4_M[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\pc_plus_4_M~3_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[2]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[2] .is_wysiwyg = "true";
defparam \pc_plus_4_M[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N21
dffeas \pc_plus_4_WB[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[2]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[2]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[2] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N5
dffeas \dmemload_WB[2] (
	.clk(CLK),
	.d(\dpif.dmemload [2]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[2]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[2] .is_wysiwyg = "true";
defparam \dmemload_WB[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N19
dffeas \porto_WB[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_2),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[2]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[2] .is_wysiwyg = "true";
defparam \porto_WB[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N18
cycloneive_lcell_comb \wdat_WB[2]~56 (
// Equation(s):
// \wdat_WB[2]~56_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[2])) # (!\memToReg_WB~q  & ((porto_WB[2])))))

	.dataa(\jal_WB~q ),
	.datab(dmemload_WB[2]),
	.datac(porto_WB[2]),
	.datad(\memToReg_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[2]~56_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[2]~56 .lut_mask = 16'h4450;
defparam \wdat_WB[2]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N20
cycloneive_lcell_comb \wdat_WB[2]~57 (
// Equation(s):
// \wdat_WB[2]~57_combout  = (!\lui_WB~q  & ((\wdat_WB[2]~56_combout ) # ((\jal_WB~q  & pc_plus_4_WB[2]))))

	.dataa(\jal_WB~q ),
	.datab(\lui_WB~q ),
	.datac(pc_plus_4_WB[2]),
	.datad(\wdat_WB[2]~56_combout ),
	.cin(gnd),
	.combout(\wdat_WB[2]~57_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[2]~57 .lut_mask = 16'h3320;
defparam \wdat_WB[2]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N4
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = (!forward_B1 & (forward_B & !Equal5))

	.dataa(\FORWARDING_UNIT|forward_B~1_combout ),
	.datab(\FORWARDING_UNIT|forward_B~0_combout ),
	.datac(gnd),
	.datad(\FORWARDING_UNIT|Equal5~1_combout ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h0044;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N4
cycloneive_lcell_comb \instruction_D~91 (
// Equation(s):
// \instruction_D~91_combout  = (iwait & (ramiframload_8 & \branch_or_jump~1_combout ))

	.dataa(iwait),
	.datab(\dpif.dmemload [8]),
	.datac(\branch_or_jump~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\instruction_D~91_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~91 .lut_mask = 16'h8080;
defparam \instruction_D~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N5
dffeas \instruction_D[8] (
	.clk(CLK),
	.d(\instruction_D~91_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[8]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[8] .is_wysiwyg = "true";
defparam \instruction_D[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N16
cycloneive_lcell_comb \imm_EX~5 (
// Equation(s):
// \imm_EX~5_combout  = (\branch_or_jump~2_combout  & (instruction_D[8] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(\branch_or_jump~2_combout ),
	.datac(\branch_taken~0_combout ),
	.datad(instruction_D[8]),
	.cin(gnd),
	.combout(\imm_EX~5_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~5 .lut_mask = 16'h8400;
defparam \imm_EX~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N17
dffeas \imm_EX[8] (
	.clk(CLK),
	.d(\imm_EX~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[8]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[8] .is_wysiwyg = "true";
defparam \imm_EX[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N6
cycloneive_lcell_comb \instruction_D~83 (
// Equation(s):
// \instruction_D~83_combout  = (\branch_or_jump~1_combout  & (ramiframload_2 & iwait))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(\dpif.dmemload [2]),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~83_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~83 .lut_mask = 16'hC000;
defparam \instruction_D~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N7
dffeas \instruction_D[2] (
	.clk(CLK),
	.d(\instruction_D~83_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[2]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[2] .is_wysiwyg = "true";
defparam \instruction_D[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N12
cycloneive_lcell_comb \instruction_D~80 (
// Equation(s):
// \instruction_D~80_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_5))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(iwait),
	.datad(ramiframload_5),
	.cin(gnd),
	.combout(\instruction_D~80_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~80 .lut_mask = 16'hA000;
defparam \instruction_D~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N13
dffeas \instruction_D[5] (
	.clk(CLK),
	.d(\instruction_D~80_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[5]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[5] .is_wysiwyg = "true";
defparam \instruction_D[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N0
cycloneive_lcell_comb \instruction_D~82 (
// Equation(s):
// \instruction_D~82_combout  = (ramiframload_3 & (\branch_or_jump~1_combout  & iwait))

	.dataa(gnd),
	.datab(ramiframload_3),
	.datac(\branch_or_jump~1_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~82_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~82 .lut_mask = 16'hC000;
defparam \instruction_D~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N1
dffeas \instruction_D[3] (
	.clk(CLK),
	.d(\instruction_D~82_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[3]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[3] .is_wysiwyg = "true";
defparam \instruction_D[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N14
cycloneive_lcell_comb \ShiftOp_EX~0 (
// Equation(s):
// \ShiftOp_EX~0_combout  = (!instruction_D[0] & (!instruction_D[2] & (!instruction_D[5] & !instruction_D[3])))

	.dataa(instruction_D[0]),
	.datab(instruction_D[2]),
	.datac(instruction_D[5]),
	.datad(instruction_D[3]),
	.cin(gnd),
	.combout(\ShiftOp_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftOp_EX~0 .lut_mask = 16'h0001;
defparam \ShiftOp_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N18
cycloneive_lcell_comb \instruction_D~85 (
// Equation(s):
// \instruction_D~85_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_4))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(ramiframload_4),
	.cin(gnd),
	.combout(\instruction_D~85_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~85 .lut_mask = 16'hC000;
defparam \instruction_D~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N19
dffeas \instruction_D[4] (
	.clk(CLK),
	.d(\instruction_D~85_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[4]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[4] .is_wysiwyg = "true";
defparam \instruction_D[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N22
cycloneive_lcell_comb \ShiftOp_EX~1 (
// Equation(s):
// \ShiftOp_EX~1_combout  = (Equal31 & (\ShiftOp_EX~0_combout  & (\branch_or_jump~1_combout  & !instruction_D[4])))

	.dataa(\CONTROL_UNIT|Equal3~2_combout ),
	.datab(\ShiftOp_EX~0_combout ),
	.datac(\branch_or_jump~1_combout ),
	.datad(instruction_D[4]),
	.cin(gnd),
	.combout(\ShiftOp_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftOp_EX~1 .lut_mask = 16'h0080;
defparam \ShiftOp_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N23
dffeas ShiftOp_EX(
	.clk(CLK),
	.d(\ShiftOp_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\ShiftOp_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam ShiftOp_EX.is_wysiwyg = "true";
defparam ShiftOp_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N26
cycloneive_lcell_comb \portB~88 (
// Equation(s):
// \portB~88_combout  = (!\Equal2~0_combout  & (!fuifforward_B_11 & ((\ALUSrc_EX~q ) # (\ShiftOp_EX~q ))))

	.dataa(\ALUSrc_EX~q ),
	.datab(\ShiftOp_EX~q ),
	.datac(\Equal2~0_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_B[1]~4_combout ),
	.cin(gnd),
	.combout(\portB~88_combout ),
	.cout());
// synopsys translate_off
defparam \portB~88 .lut_mask = 16'h000E;
defparam \portB~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N8
cycloneive_lcell_comb \portB~93 (
// Equation(s):
// \portB~93_combout  = (\ShiftOp_EX~q ) # ((\Equal2~0_combout ) # (fuifforward_B_11))

	.dataa(gnd),
	.datab(\ShiftOp_EX~q ),
	.datac(\Equal2~0_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_B[1]~4_combout ),
	.cin(gnd),
	.combout(\portB~93_combout ),
	.cout());
// synopsys translate_off
defparam \portB~93 .lut_mask = 16'hFFFC;
defparam \portB~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N6
cycloneive_lcell_comb \portB~98 (
// Equation(s):
// \portB~98_combout  = (\portB~88_combout  & (((\portB~93_combout )))) # (!\portB~88_combout  & ((\portB~93_combout  & ((\wdat_WB[2]~57_combout ))) # (!\portB~93_combout  & (rdata2_EX[2]))))

	.dataa(rdata2_EX[2]),
	.datab(\wdat_WB[2]~57_combout ),
	.datac(\portB~88_combout ),
	.datad(\portB~93_combout ),
	.cin(gnd),
	.combout(\portB~98_combout ),
	.cout());
// synopsys translate_off
defparam \portB~98 .lut_mask = 16'hFC0A;
defparam \portB~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N24
cycloneive_lcell_comb \portB~99 (
// Equation(s):
// \portB~99_combout  = (\portB~88_combout  & ((\portB~98_combout  & ((imm_EX[8]))) # (!\portB~98_combout  & (imm_EX[2])))) # (!\portB~88_combout  & (((\portB~98_combout ))))

	.dataa(imm_EX[2]),
	.datab(imm_EX[8]),
	.datac(\portB~88_combout ),
	.datad(\portB~98_combout ),
	.cin(gnd),
	.combout(\portB~99_combout ),
	.cout());
// synopsys translate_off
defparam \portB~99 .lut_mask = 16'hCFA0;
defparam \portB~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N30
cycloneive_lcell_comb \portB~100 (
// Equation(s):
// \portB~100_combout  = (\Equal2~0_combout  & (porto_M_2 & (!\lui_M~q ))) # (!\Equal2~0_combout  & (((\portB~99_combout ))))

	.dataa(porto_M_2),
	.datab(\lui_M~q ),
	.datac(\Equal2~0_combout ),
	.datad(\portB~99_combout ),
	.cin(gnd),
	.combout(\portB~100_combout ),
	.cout());
// synopsys translate_off
defparam \portB~100 .lut_mask = 16'h2F20;
defparam \portB~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N18
cycloneive_lcell_comb \rdata2_EX~58 (
// Equation(s):
// \rdata2_EX~58_combout  = (instruction_D[20] & (Mux61)) # (!instruction_D[20] & ((Mux611)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux61~9_combout ),
	.datad(\REGISTER_FILE|Mux61~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~58_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~58 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N18
cycloneive_lcell_comb \rdata2_EX~59 (
// Equation(s):
// \rdata2_EX~59_combout  = (\always2~2_combout  & ((\rdata2_EX~58_combout ))) # (!\always2~2_combout  & (\portB~100_combout ))

	.dataa(\always2~2_combout ),
	.datab(gnd),
	.datac(\portB~100_combout ),
	.datad(\rdata2_EX~58_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~59_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~59 .lut_mask = 16'hFA50;
defparam \rdata2_EX~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N30
cycloneive_lcell_comb \Equal3~2 (
// Equation(s):
// \Equal3~2_combout  = (fuifforward_B_11) # ((!forward_B1 & (!Equal5 & forward_B)))

	.dataa(\FORWARDING_UNIT|forward_B~1_combout ),
	.datab(\FORWARDING_UNIT|Equal5~1_combout ),
	.datac(\FORWARDING_UNIT|forward_B~0_combout ),
	.datad(\FORWARDING_UNIT|fuif.forward_B[1]~4_combout ),
	.cin(gnd),
	.combout(\Equal3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~2 .lut_mask = 16'hFF10;
defparam \Equal3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N6
cycloneive_lcell_comb \rdata1_EX[15]~0 (
// Equation(s):
// \rdata1_EX[15]~0_combout  = ((!fuifforward_A_01 & (!\Equal3~2_combout  & !fuifforward_A_11))) # (!dREN_M1)

	.dataa(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datab(\Equal3~2_combout ),
	.datac(dREN_M1),
	.datad(\FORWARDING_UNIT|fuif.forward_A[1]~7_combout ),
	.cin(gnd),
	.combout(\rdata1_EX[15]~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX[15]~0 .lut_mask = 16'h0F1F;
defparam \rdata1_EX[15]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N20
cycloneive_lcell_comb \always2~2 (
// Equation(s):
// \always2~2_combout  = (((!dREN_M1 & !dWEN_M1)) # (!fuifbubble_lw_f)) # (!always1)

	.dataa(dREN_M1),
	.datab(dWEN_M1),
	.datac(always1),
	.datad(\FORWARDING_UNIT|fuif.bubble_lw_f~2_combout ),
	.cin(gnd),
	.combout(\always2~2_combout ),
	.cout());
// synopsys translate_off
defparam \always2~2 .lut_mask = 16'h1FFF;
defparam \always2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N26
cycloneive_lcell_comb \rdata1_EX[15]~1 (
// Equation(s):
// \rdata1_EX[15]~1_combout  = ((!\en_EX~0_combout  & ((\always2~2_combout ) # (!\rdata1_EX[15]~0_combout )))) # (!\branch_or_jump~1_combout )

	.dataa(\branch_or_jump~1_combout ),
	.datab(\rdata1_EX[15]~0_combout ),
	.datac(\en_EX~0_combout ),
	.datad(\always2~2_combout ),
	.cin(gnd),
	.combout(\rdata1_EX[15]~1_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX[15]~1 .lut_mask = 16'h5F57;
defparam \rdata1_EX[15]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N19
dffeas \rdata2_EX[2] (
	.clk(CLK),
	.d(\rdata2_EX~59_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[2]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[2] .is_wysiwyg = "true";
defparam \rdata2_EX[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N6
cycloneive_lcell_comb \rdata2_M~6 (
// Equation(s):
// \rdata2_M~6_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & ((\rdata2_M[16]~1_combout  & (\sw_forwarding_output~29_combout )) # (!\rdata2_M[16]~1_combout  & ((rdata2_EX[2])))))

	.dataa(\sw_forwarding_output~29_combout ),
	.datab(rdata2_EX[2]),
	.datac(\rdata2_M[16]~0_combout ),
	.datad(\rdata2_M[16]~1_combout ),
	.cin(gnd),
	.combout(\rdata2_M~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~6 .lut_mask = 16'hFA0C;
defparam \rdata2_M~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N24
cycloneive_lcell_comb \rdata2_M~7 (
// Equation(s):
// \rdata2_M~7_combout  = (\rdata2_M[16]~0_combout  & ((\rdata2_M~6_combout  & (\wdat_WB[2]~57_combout )) # (!\rdata2_M~6_combout  & ((ramiframload_2))))) # (!\rdata2_M[16]~0_combout  & (((\rdata2_M~6_combout ))))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(\wdat_WB[2]~57_combout ),
	.datac(\dpif.dmemload [2]),
	.datad(\rdata2_M~6_combout ),
	.cin(gnd),
	.combout(\rdata2_M~7_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~7 .lut_mask = 16'hDDA0;
defparam \rdata2_M~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N28
cycloneive_lcell_comb \pc_plus_4_EX~2 (
// Equation(s):
// \pc_plus_4_EX~2_combout  = (pc_plus_4_D[3] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[3]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~2 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N29
dffeas \pc_plus_4_EX[3] (
	.clk(CLK),
	.d(\pc_plus_4_EX~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[3]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[3] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N12
cycloneive_lcell_comb \pc_plus_4_M~2 (
// Equation(s):
// \pc_plus_4_M~2_combout  = (pc_plus_4_EX[3] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[3]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~2_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~2 .lut_mask = 16'h00CC;
defparam \pc_plus_4_M~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N13
dffeas \pc_plus_4_M[3] (
	.clk(CLK),
	.d(\pc_plus_4_M~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[3]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[3] .is_wysiwyg = "true";
defparam \pc_plus_4_M[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N3
dffeas \pc_plus_4_WB[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[3]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[3]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[3] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N1
dffeas \porto_WB[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_3),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[3]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[3] .is_wysiwyg = "true";
defparam \porto_WB[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N0
cycloneive_lcell_comb \wdat_WB[3]~64 (
// Equation(s):
// \wdat_WB[3]~64_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[3])) # (!\memToReg_WB~q  & ((porto_WB[3])))))

	.dataa(dmemload_WB[3]),
	.datab(\jal_WB~q ),
	.datac(porto_WB[3]),
	.datad(\memToReg_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[3]~64_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[3]~64 .lut_mask = 16'h2230;
defparam \wdat_WB[3]~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N2
cycloneive_lcell_comb \wdat_WB[3]~65 (
// Equation(s):
// \wdat_WB[3]~65_combout  = (!\lui_WB~q  & ((\wdat_WB[3]~64_combout ) # ((\jal_WB~q  & pc_plus_4_WB[3]))))

	.dataa(\lui_WB~q ),
	.datab(\jal_WB~q ),
	.datac(pc_plus_4_WB[3]),
	.datad(\wdat_WB[3]~64_combout ),
	.cin(gnd),
	.combout(\wdat_WB[3]~65_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[3]~65 .lut_mask = 16'h5540;
defparam \wdat_WB[3]~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N14
cycloneive_lcell_comb \rdata2_M~8 (
// Equation(s):
// \rdata2_M~8_combout  = (\rdata2_M[16]~1_combout  & (((\rdata2_M[16]~0_combout )))) # (!\rdata2_M[16]~1_combout  & ((\rdata2_M[16]~0_combout  & ((ramiframload_3))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[3]))))

	.dataa(rdata2_EX[3]),
	.datab(\rdata2_M[16]~1_combout ),
	.datac(ramiframload_3),
	.datad(\rdata2_M[16]~0_combout ),
	.cin(gnd),
	.combout(\rdata2_M~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~8 .lut_mask = 16'hFC22;
defparam \rdata2_M~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N22
cycloneive_lcell_comb \sw_forwarding_output~30 (
// Equation(s):
// \sw_forwarding_output~30_combout  = (!\lui_M~q  & porto_M_3)

	.dataa(gnd),
	.datab(\lui_M~q ),
	.datac(gnd),
	.datad(porto_M_3),
	.cin(gnd),
	.combout(\sw_forwarding_output~30_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~30 .lut_mask = 16'h3300;
defparam \sw_forwarding_output~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N0
cycloneive_lcell_comb \rdata2_M~9 (
// Equation(s):
// \rdata2_M~9_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~8_combout  & (\wdat_WB[3]~65_combout )) # (!\rdata2_M~8_combout  & ((\sw_forwarding_output~30_combout ))))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~8_combout ))))

	.dataa(\wdat_WB[3]~65_combout ),
	.datab(\rdata2_M[16]~1_combout ),
	.datac(\rdata2_M~8_combout ),
	.datad(\sw_forwarding_output~30_combout ),
	.cin(gnd),
	.combout(\rdata2_M~9_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~9 .lut_mask = 16'hBCB0;
defparam \rdata2_M~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N26
cycloneive_lcell_comb \portB~104 (
// Equation(s):
// \portB~104_combout  = (\portB~93_combout  & (\wdat_WB[4]~63_combout )) # (!\portB~93_combout  & ((rdata2_EX[4])))

	.dataa(\wdat_WB[4]~63_combout ),
	.datab(rdata2_EX[4]),
	.datac(\portB~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\portB~104_combout ),
	.cout());
// synopsys translate_off
defparam \portB~104 .lut_mask = 16'hACAC;
defparam \portB~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N18
cycloneive_lcell_comb \imm_EX~15 (
// Equation(s):
// \imm_EX~15_combout  = (instruction_D[4] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(\branch_taken~0_combout ),
	.datac(instruction_D[4]),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\imm_EX~15_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~15 .lut_mask = 16'h9000;
defparam \imm_EX~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N19
dffeas \imm_EX[4] (
	.clk(CLK),
	.d(\imm_EX~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[4]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[4] .is_wysiwyg = "true";
defparam \imm_EX[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N4
cycloneive_lcell_comb \portB~105 (
// Equation(s):
// \portB~105_combout  = (\Equal2~0_combout  & (porto_M_4 & (!\lui_M~q ))) # (!\Equal2~0_combout  & (((imm_EX[4]))))

	.dataa(porto_M_4),
	.datab(\lui_M~q ),
	.datac(\Equal2~0_combout ),
	.datad(imm_EX[4]),
	.cin(gnd),
	.combout(\portB~105_combout ),
	.cout());
// synopsys translate_off
defparam \portB~105 .lut_mask = 16'h2F20;
defparam \portB~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N16
cycloneive_lcell_comb \instruction_D~93 (
// Equation(s):
// \instruction_D~93_combout  = (ramiframload_10 & (\branch_or_jump~1_combout  & iwait))

	.dataa(gnd),
	.datab(\dpif.dmemload [10]),
	.datac(\branch_or_jump~1_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~93_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~93 .lut_mask = 16'hC000;
defparam \instruction_D~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N17
dffeas \instruction_D[10] (
	.clk(CLK),
	.d(\instruction_D~93_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[10]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[10] .is_wysiwyg = "true";
defparam \instruction_D[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N28
cycloneive_lcell_comb \imm_EX~7 (
// Equation(s):
// \imm_EX~7_combout  = (\branch_or_jump~2_combout  & (instruction_D[10] & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_taken~0_combout ),
	.datab(\predicted_M~q ),
	.datac(\branch_or_jump~2_combout ),
	.datad(instruction_D[10]),
	.cin(gnd),
	.combout(\imm_EX~7_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~7 .lut_mask = 16'h9000;
defparam \imm_EX~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N29
dffeas \imm_EX[10] (
	.clk(CLK),
	.d(\imm_EX~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[10]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[10] .is_wysiwyg = "true";
defparam \imm_EX[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N6
cycloneive_lcell_comb \portB~106 (
// Equation(s):
// \portB~106_combout  = (\Equal2~0_combout  & (\portB~105_combout )) # (!\Equal2~0_combout  & ((\portB~93_combout  & ((imm_EX[10]))) # (!\portB~93_combout  & (\portB~105_combout ))))

	.dataa(\Equal2~0_combout ),
	.datab(\portB~105_combout ),
	.datac(\portB~93_combout ),
	.datad(imm_EX[10]),
	.cin(gnd),
	.combout(\portB~106_combout ),
	.cout());
// synopsys translate_off
defparam \portB~106 .lut_mask = 16'hDC8C;
defparam \portB~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N8
cycloneive_lcell_comb \portB~107 (
// Equation(s):
// \portB~107_combout  = (\portB~88_combout  & (((\portB~106_combout )))) # (!\portB~88_combout  & ((\Equal2~0_combout  & ((\portB~106_combout ))) # (!\Equal2~0_combout  & (\portB~104_combout ))))

	.dataa(\portB~88_combout ),
	.datab(\Equal2~0_combout ),
	.datac(\portB~104_combout ),
	.datad(\portB~106_combout ),
	.cin(gnd),
	.combout(\portB~107_combout ),
	.cout());
// synopsys translate_off
defparam \portB~107 .lut_mask = 16'hFE10;
defparam \portB~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N4
cycloneive_lcell_comb \instruction_D~74 (
// Equation(s):
// \instruction_D~74_combout  = (\branch_or_jump~1_combout  & (ramiframload_20 & iwait))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(ramiframload_20),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~74_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~74 .lut_mask = 16'hC000;
defparam \instruction_D~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N5
dffeas \instruction_D[20] (
	.clk(CLK),
	.d(\instruction_D~74_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[20]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[20] .is_wysiwyg = "true";
defparam \instruction_D[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N20
cycloneive_lcell_comb \rdata2_EX~62 (
// Equation(s):
// \rdata2_EX~62_combout  = (instruction_D[20] & ((Mux59))) # (!instruction_D[20] & (Mux591))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux59~19_combout ),
	.datad(\REGISTER_FILE|Mux59~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~62_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~62 .lut_mask = 16'hFC30;
defparam \rdata2_EX~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N14
cycloneive_lcell_comb \rdata2_EX~63 (
// Equation(s):
// \rdata2_EX~63_combout  = (\always2~2_combout  & ((\rdata2_EX~62_combout ))) # (!\always2~2_combout  & (\portB~107_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portB~107_combout ),
	.datad(\rdata2_EX~62_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~63_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~63 .lut_mask = 16'hFC30;
defparam \rdata2_EX~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N15
dffeas \rdata2_EX[4] (
	.clk(CLK),
	.d(\rdata2_EX~63_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[4]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[4] .is_wysiwyg = "true";
defparam \rdata2_EX[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N10
cycloneive_lcell_comb \rdata2_M~10 (
// Equation(s):
// \rdata2_M~10_combout  = (\rdata2_M[16]~1_combout  & ((\sw_forwarding_output~31_combout ) # ((\rdata2_M[16]~0_combout )))) # (!\rdata2_M[16]~1_combout  & (((rdata2_EX[4] & !\rdata2_M[16]~0_combout ))))

	.dataa(\sw_forwarding_output~31_combout ),
	.datab(rdata2_EX[4]),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\rdata2_M[16]~0_combout ),
	.cin(gnd),
	.combout(\rdata2_M~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~10 .lut_mask = 16'hF0AC;
defparam \rdata2_M~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N2
cycloneive_lcell_comb \pc_plus_4_EX~5 (
// Equation(s):
// \pc_plus_4_EX~5_combout  = (pc_plus_4_D[4] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[4]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~5_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~5 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N3
dffeas \pc_plus_4_EX[4] (
	.clk(CLK),
	.d(\pc_plus_4_EX~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[4]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[4] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N18
cycloneive_lcell_comb \pc_plus_4_M~5 (
// Equation(s):
// \pc_plus_4_M~5_combout  = (pc_plus_4_EX[4] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[4]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~5_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~5 .lut_mask = 16'h00CC;
defparam \pc_plus_4_M~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N19
dffeas \pc_plus_4_M[4] (
	.clk(CLK),
	.d(\pc_plus_4_M~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[4]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[4] .is_wysiwyg = "true";
defparam \pc_plus_4_M[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N29
dffeas \pc_plus_4_WB[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[4]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[4]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[4] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N28
cycloneive_lcell_comb \wdat_WB[4]~63 (
// Equation(s):
// \wdat_WB[4]~63_combout  = (!\lui_WB~q  & ((\wdat_WB[4]~62_combout ) # ((\jal_WB~q  & pc_plus_4_WB[4]))))

	.dataa(\wdat_WB[4]~62_combout ),
	.datab(\jal_WB~q ),
	.datac(pc_plus_4_WB[4]),
	.datad(\lui_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[4]~63_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[4]~63 .lut_mask = 16'h00EA;
defparam \wdat_WB[4]~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N20
cycloneive_lcell_comb \rdata2_M~11 (
// Equation(s):
// \rdata2_M~11_combout  = (\rdata2_M~10_combout  & (((\wdat_WB[4]~63_combout )) # (!\rdata2_M[16]~0_combout ))) # (!\rdata2_M~10_combout  & (\rdata2_M[16]~0_combout  & ((ramiframload_4))))

	.dataa(\rdata2_M~10_combout ),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\wdat_WB[4]~63_combout ),
	.datad(ramiframload_4),
	.cin(gnd),
	.combout(\rdata2_M~11_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~11 .lut_mask = 16'hE6A2;
defparam \rdata2_M~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N28
cycloneive_lcell_comb \pc_plus_4_EX~4 (
// Equation(s):
// \pc_plus_4_EX~4_combout  = (pc_plus_4_D[5] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[5]),
	.datab(\predicted_M~q ),
	.datac(\branch_or_jump~2_combout ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~4_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~4 .lut_mask = 16'h8020;
defparam \pc_plus_4_EX~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N29
dffeas \pc_plus_4_EX[5] (
	.clk(CLK),
	.d(\pc_plus_4_EX~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[5]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[5] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N10
cycloneive_lcell_comb \pc_plus_4_M~4 (
// Equation(s):
// \pc_plus_4_M~4_combout  = (pc_plus_4_EX[5] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_plus_4_EX[5]),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~4_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~4 .lut_mask = 16'h00F0;
defparam \pc_plus_4_M~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N11
dffeas \pc_plus_4_M[5] (
	.clk(CLK),
	.d(\pc_plus_4_M~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[5]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[5] .is_wysiwyg = "true";
defparam \pc_plus_4_M[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N15
dffeas \pc_plus_4_WB[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[5]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[5]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[5] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N23
dffeas \dmemload_WB[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_5),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[5]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[5] .is_wysiwyg = "true";
defparam \dmemload_WB[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N17
dffeas \porto_WB[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_5),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[5]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[5] .is_wysiwyg = "true";
defparam \porto_WB[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N16
cycloneive_lcell_comb \wdat_WB[5]~54 (
// Equation(s):
// \wdat_WB[5]~54_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[5])) # (!\memToReg_WB~q  & ((porto_WB[5])))))

	.dataa(\memToReg_WB~q ),
	.datab(dmemload_WB[5]),
	.datac(porto_WB[5]),
	.datad(\jal_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[5]~54_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[5]~54 .lut_mask = 16'h00D8;
defparam \wdat_WB[5]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N14
cycloneive_lcell_comb \wdat_WB[5]~55 (
// Equation(s):
// \wdat_WB[5]~55_combout  = (!\lui_WB~q  & ((\wdat_WB[5]~54_combout ) # ((\jal_WB~q  & pc_plus_4_WB[5]))))

	.dataa(\jal_WB~q ),
	.datab(\lui_WB~q ),
	.datac(pc_plus_4_WB[5]),
	.datad(\wdat_WB[5]~54_combout ),
	.cin(gnd),
	.combout(\wdat_WB[5]~55_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[5]~55 .lut_mask = 16'h3320;
defparam \wdat_WB[5]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N16
cycloneive_lcell_comb \sw_forwarding_output~26 (
// Equation(s):
// \sw_forwarding_output~26_combout  = (!\lui_M~q  & porto_M_5)

	.dataa(\lui_M~q ),
	.datab(gnd),
	.datac(porto_M_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\sw_forwarding_output~26_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~26 .lut_mask = 16'h5050;
defparam \sw_forwarding_output~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N10
cycloneive_lcell_comb \rdata2_M~12 (
// Equation(s):
// \rdata2_M~12_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout ) # (ramiframload_5)))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[5] & (!\rdata2_M[16]~1_combout )))

	.dataa(rdata2_EX[5]),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(ramiframload_5),
	.cin(gnd),
	.combout(\rdata2_M~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~12 .lut_mask = 16'hCEC2;
defparam \rdata2_M~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N0
cycloneive_lcell_comb \rdata2_M~13 (
// Equation(s):
// \rdata2_M~13_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~12_combout  & (\wdat_WB[5]~55_combout )) # (!\rdata2_M~12_combout  & ((\sw_forwarding_output~26_combout ))))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~12_combout ))))

	.dataa(\wdat_WB[5]~55_combout ),
	.datab(\sw_forwarding_output~26_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\rdata2_M~12_combout ),
	.cin(gnd),
	.combout(\rdata2_M~13_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~13 .lut_mask = 16'hAFC0;
defparam \rdata2_M~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N8
cycloneive_lcell_comb \pc_plus_4_EX~7 (
// Equation(s):
// \pc_plus_4_EX~7_combout  = (pc_plus_4_D[6] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(pc_plus_4_D[6]),
	.datab(\branch_taken~0_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~7_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~7 .lut_mask = 16'h8200;
defparam \pc_plus_4_EX~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N9
dffeas \pc_plus_4_EX[6] (
	.clk(CLK),
	.d(\pc_plus_4_EX~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[6]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[6] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N14
cycloneive_lcell_comb \pc_plus_4_M~7 (
// Equation(s):
// \pc_plus_4_M~7_combout  = (pc_plus_4_EX[6] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_plus_4_EX[6]),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~7_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~7 .lut_mask = 16'h00F0;
defparam \pc_plus_4_M~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y36_N15
dffeas \pc_plus_4_M[6] (
	.clk(CLK),
	.d(\pc_plus_4_M~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[6]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[6] .is_wysiwyg = "true";
defparam \pc_plus_4_M[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N7
dffeas \pc_plus_4_WB[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[6]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[6]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[6] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N9
dffeas \porto_WB[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_6),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[6]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[6] .is_wysiwyg = "true";
defparam \porto_WB[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N8
cycloneive_lcell_comb \wdat_WB[6]~52 (
// Equation(s):
// \wdat_WB[6]~52_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[6])) # (!\memToReg_WB~q  & ((porto_WB[6])))))

	.dataa(dmemload_WB[6]),
	.datab(\jal_WB~q ),
	.datac(porto_WB[6]),
	.datad(\memToReg_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[6]~52_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[6]~52 .lut_mask = 16'h2230;
defparam \wdat_WB[6]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N6
cycloneive_lcell_comb \wdat_WB[6]~53 (
// Equation(s):
// \wdat_WB[6]~53_combout  = (!\lui_WB~q  & ((\wdat_WB[6]~52_combout ) # ((\jal_WB~q  & pc_plus_4_WB[6]))))

	.dataa(\lui_WB~q ),
	.datab(\jal_WB~q ),
	.datac(pc_plus_4_WB[6]),
	.datad(\wdat_WB[6]~52_combout ),
	.cin(gnd),
	.combout(\wdat_WB[6]~53_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[6]~53 .lut_mask = 16'h5540;
defparam \wdat_WB[6]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N4
cycloneive_lcell_comb \instruction_D~95 (
// Equation(s):
// \instruction_D~95_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_6))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(\dpif.dmemload [6]),
	.cin(gnd),
	.combout(\instruction_D~95_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~95 .lut_mask = 16'hC000;
defparam \instruction_D~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N5
dffeas \instruction_D[6] (
	.clk(CLK),
	.d(\instruction_D~95_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[6]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[6] .is_wysiwyg = "true";
defparam \instruction_D[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N18
cycloneive_lcell_comb \imm_EX~9 (
// Equation(s):
// \imm_EX~9_combout  = (instruction_D[6] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_taken~0_combout ),
	.datab(instruction_D[6]),
	.datac(\predicted_M~q ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\imm_EX~9_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~9 .lut_mask = 16'h8400;
defparam \imm_EX~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N29
dffeas \imm_EX[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\imm_EX~9_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[6]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[6] .is_wysiwyg = "true";
defparam \imm_EX[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N20
cycloneive_lcell_comb \portB~14 (
// Equation(s):
// \portB~14_combout  = (\Equal2~0_combout ) # ((\ALUSrc_EX~q  & !fuifforward_B_11))

	.dataa(\ALUSrc_EX~q ),
	.datab(\Equal2~0_combout ),
	.datac(gnd),
	.datad(\FORWARDING_UNIT|fuif.forward_B[1]~4_combout ),
	.cin(gnd),
	.combout(\portB~14_combout ),
	.cout());
// synopsys translate_off
defparam \portB~14 .lut_mask = 16'hCCEE;
defparam \portB~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N0
cycloneive_lcell_comb \portB~83 (
// Equation(s):
// \portB~83_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & (imm_EX[6])) # (!\portB~14_combout  & ((rdata2_EX[6])))))

	.dataa(\ShiftOp_EX~q ),
	.datab(imm_EX[6]),
	.datac(rdata2_EX[6]),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~83_combout ),
	.cout());
// synopsys translate_off
defparam \portB~83 .lut_mask = 16'h4450;
defparam \portB~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N10
cycloneive_lcell_comb \portB~115 (
// Equation(s):
// \portB~115_combout  = (\portB~14_combout  & (porto_M_6 & ((!\lui_M~q )))) # (!\portB~14_combout  & (((\wdat_WB[6]~53_combout ))))

	.dataa(porto_M_6),
	.datab(\wdat_WB[6]~53_combout ),
	.datac(\lui_M~q ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~115_combout ),
	.cout());
// synopsys translate_off
defparam \portB~115 .lut_mask = 16'h0ACC;
defparam \portB~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N20
cycloneive_lcell_comb \portB~84 (
// Equation(s):
// \portB~84_combout  = (\Equal3~2_combout  & ((\portB~115_combout ))) # (!\Equal3~2_combout  & (\portB~83_combout ))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~83_combout ),
	.datad(\portB~115_combout ),
	.cin(gnd),
	.combout(\portB~84_combout ),
	.cout());
// synopsys translate_off
defparam \portB~84 .lut_mask = 16'hFA50;
defparam \portB~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N12
cycloneive_lcell_comb \rdata2_EX~50 (
// Equation(s):
// \rdata2_EX~50_combout  = (instruction_D[20] & ((Mux57))) # (!instruction_D[20] & (Mux571))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux57~19_combout ),
	.datad(\REGISTER_FILE|Mux57~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~50_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~50 .lut_mask = 16'hFA50;
defparam \rdata2_EX~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N4
cycloneive_lcell_comb \rdata2_EX~51 (
// Equation(s):
// \rdata2_EX~51_combout  = (\always2~2_combout  & ((\rdata2_EX~50_combout ))) # (!\always2~2_combout  & (\portB~84_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portB~84_combout ),
	.datad(\rdata2_EX~50_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~51_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~51 .lut_mask = 16'hFC30;
defparam \rdata2_EX~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N5
dffeas \rdata2_EX[6] (
	.clk(CLK),
	.d(\rdata2_EX~51_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[6]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[6] .is_wysiwyg = "true";
defparam \rdata2_EX[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N8
cycloneive_lcell_comb \rdata2_M~14 (
// Equation(s):
// \rdata2_M~14_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & ((\rdata2_M[16]~1_combout  & (\sw_forwarding_output~25_combout )) # (!\rdata2_M[16]~1_combout  & ((rdata2_EX[6])))))

	.dataa(\sw_forwarding_output~25_combout ),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(rdata2_EX[6]),
	.datad(\rdata2_M[16]~1_combout ),
	.cin(gnd),
	.combout(\rdata2_M~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~14 .lut_mask = 16'hEE30;
defparam \rdata2_M~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N10
cycloneive_lcell_comb \rdata2_M~15 (
// Equation(s):
// \rdata2_M~15_combout  = (\rdata2_M[16]~0_combout  & ((\rdata2_M~14_combout  & (\wdat_WB[6]~53_combout )) # (!\rdata2_M~14_combout  & ((ramiframload_6))))) # (!\rdata2_M[16]~0_combout  & (((\rdata2_M~14_combout ))))

	.dataa(\wdat_WB[6]~53_combout ),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\rdata2_M~14_combout ),
	.datad(\dpif.dmemload [6]),
	.cin(gnd),
	.combout(\rdata2_M~15_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~15 .lut_mask = 16'hBCB0;
defparam \rdata2_M~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N26
cycloneive_lcell_comb \sw_forwarding_output~24 (
// Equation(s):
// \sw_forwarding_output~24_combout  = (!\lui_M~q  & porto_M_7)

	.dataa(\lui_M~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(porto_M_7),
	.cin(gnd),
	.combout(\sw_forwarding_output~24_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~24 .lut_mask = 16'h5500;
defparam \sw_forwarding_output~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N12
cycloneive_lcell_comb \pc_plus_4[7]~10 (
// Equation(s):
// \pc_plus_4[7]~10_combout  = (pc_out_7 & (!\pc_plus_4[6]~9 )) # (!pc_out_7 & ((\pc_plus_4[6]~9 ) # (GND)))
// \pc_plus_4[7]~11  = CARRY((!\pc_plus_4[6]~9 ) # (!pc_out_7))

	.dataa(pc_out_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[6]~9 ),
	.combout(\pc_plus_4[7]~10_combout ),
	.cout(\pc_plus_4[7]~11 ));
// synopsys translate_off
defparam \pc_plus_4[7]~10 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[7]~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N16
cycloneive_lcell_comb \pc_plus_4_D~6 (
// Equation(s):
// \pc_plus_4_D~6_combout  = (\pc_plus_4[7]~10_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(\pc_plus_4[7]~10_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\pc_plus_4_D~6_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~6 .lut_mask = 16'hF050;
defparam \pc_plus_4_D~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N17
dffeas \pc_plus_4_D[7] (
	.clk(CLK),
	.d(\pc_plus_4_D~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[7]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[7] .is_wysiwyg = "true";
defparam \pc_plus_4_D[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N24
cycloneive_lcell_comb \pc_plus_4_EX~6 (
// Equation(s):
// \pc_plus_4_EX~6_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[7] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_D[7]),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~6_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~6 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N25
dffeas \pc_plus_4_EX[7] (
	.clk(CLK),
	.d(\pc_plus_4_EX~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[7]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[7] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N8
cycloneive_lcell_comb \pc_plus_4_M~6 (
// Equation(s):
// \pc_plus_4_M~6_combout  = (pc_plus_4_EX[7] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[7]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~6_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~6 .lut_mask = 16'h00CC;
defparam \pc_plus_4_M~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N9
dffeas \pc_plus_4_M[7] (
	.clk(CLK),
	.d(\pc_plus_4_M~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[7]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[7] .is_wysiwyg = "true";
defparam \pc_plus_4_M[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N13
dffeas \pc_plus_4_WB[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[7]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[7]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[7] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N4
cycloneive_lcell_comb \dmemload_WB[7]~feeder (
// Equation(s):
// \dmemload_WB[7]~feeder_combout  = ramiframload_7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_7),
	.cin(gnd),
	.combout(\dmemload_WB[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \dmemload_WB[7]~feeder .lut_mask = 16'hFF00;
defparam \dmemload_WB[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N5
dffeas \dmemload_WB[7] (
	.clk(CLK),
	.d(\dmemload_WB[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[7]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[7] .is_wysiwyg = "true";
defparam \dmemload_WB[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N11
dffeas \porto_WB[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_7),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[7]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[7] .is_wysiwyg = "true";
defparam \porto_WB[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N10
cycloneive_lcell_comb \wdat_WB[7]~50 (
// Equation(s):
// \wdat_WB[7]~50_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[7])) # (!\memToReg_WB~q  & ((porto_WB[7])))))

	.dataa(\jal_WB~q ),
	.datab(dmemload_WB[7]),
	.datac(porto_WB[7]),
	.datad(\memToReg_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[7]~50_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[7]~50 .lut_mask = 16'h4450;
defparam \wdat_WB[7]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N12
cycloneive_lcell_comb \wdat_WB[7]~51 (
// Equation(s):
// \wdat_WB[7]~51_combout  = (!\lui_WB~q  & ((\wdat_WB[7]~50_combout ) # ((\jal_WB~q  & pc_plus_4_WB[7]))))

	.dataa(\lui_WB~q ),
	.datab(\jal_WB~q ),
	.datac(pc_plus_4_WB[7]),
	.datad(\wdat_WB[7]~50_combout ),
	.cin(gnd),
	.combout(\wdat_WB[7]~51_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[7]~51 .lut_mask = 16'h5540;
defparam \wdat_WB[7]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N28
cycloneive_lcell_comb \rdata2_M~16 (
// Equation(s):
// \rdata2_M~16_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout ) # (ramiframload_7)))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[7] & (!\rdata2_M[16]~1_combout )))

	.dataa(rdata2_EX[7]),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(ramiframload_7),
	.cin(gnd),
	.combout(\rdata2_M~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~16 .lut_mask = 16'hCEC2;
defparam \rdata2_M~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N14
cycloneive_lcell_comb \rdata2_M~17 (
// Equation(s):
// \rdata2_M~17_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~16_combout  & ((\wdat_WB[7]~51_combout ))) # (!\rdata2_M~16_combout  & (\sw_forwarding_output~24_combout )))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~16_combout ))))

	.dataa(\sw_forwarding_output~24_combout ),
	.datab(\wdat_WB[7]~51_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\rdata2_M~16_combout ),
	.cin(gnd),
	.combout(\rdata2_M~17_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~17 .lut_mask = 16'hCFA0;
defparam \rdata2_M~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N16
cycloneive_lcell_comb \pc_plus_4_M~9 (
// Equation(s):
// \pc_plus_4_M~9_combout  = (pc_plus_4_EX[8] & !\wsel_M~0_combout )

	.dataa(pc_plus_4_EX[8]),
	.datab(gnd),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~9_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~9 .lut_mask = 16'h00AA;
defparam \pc_plus_4_M~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N17
dffeas \pc_plus_4_M[8] (
	.clk(CLK),
	.d(\pc_plus_4_M~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[8]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[8] .is_wysiwyg = "true";
defparam \pc_plus_4_M[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N31
dffeas \pc_plus_4_WB[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[8]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[8]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[8] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N17
dffeas \porto_WB[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_8),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[8]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[8] .is_wysiwyg = "true";
defparam \porto_WB[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N16
cycloneive_lcell_comb \wdat_WB[8]~44 (
// Equation(s):
// \wdat_WB[8]~44_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[8])) # (!\memToReg_WB~q  & ((porto_WB[8])))))

	.dataa(dmemload_WB[8]),
	.datab(\jal_WB~q ),
	.datac(porto_WB[8]),
	.datad(\memToReg_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[8]~44_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[8]~44 .lut_mask = 16'h2230;
defparam \wdat_WB[8]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N30
cycloneive_lcell_comb \wdat_WB[8]~45 (
// Equation(s):
// \wdat_WB[8]~45_combout  = (!\lui_WB~q  & ((\wdat_WB[8]~44_combout ) # ((\jal_WB~q  & pc_plus_4_WB[8]))))

	.dataa(\lui_WB~q ),
	.datab(\jal_WB~q ),
	.datac(pc_plus_4_WB[8]),
	.datad(\wdat_WB[8]~44_combout ),
	.cin(gnd),
	.combout(\wdat_WB[8]~45_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[8]~45 .lut_mask = 16'h5540;
defparam \wdat_WB[8]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N6
cycloneive_lcell_comb \sw_forwarding_output~21 (
// Equation(s):
// \sw_forwarding_output~21_combout  = (porto_M_8 & !\lui_M~q )

	.dataa(gnd),
	.datab(gnd),
	.datac(porto_M_8),
	.datad(\lui_M~q ),
	.cin(gnd),
	.combout(\sw_forwarding_output~21_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~21 .lut_mask = 16'h00F0;
defparam \sw_forwarding_output~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N8
cycloneive_lcell_comb \rdata2_M~18 (
// Equation(s):
// \rdata2_M~18_combout  = (\rdata2_M[16]~1_combout  & (((\rdata2_M[16]~0_combout ) # (\sw_forwarding_output~21_combout )))) # (!\rdata2_M[16]~1_combout  & (rdata2_EX[8] & (!\rdata2_M[16]~0_combout )))

	.dataa(rdata2_EX[8]),
	.datab(\rdata2_M[16]~1_combout ),
	.datac(\rdata2_M[16]~0_combout ),
	.datad(\sw_forwarding_output~21_combout ),
	.cin(gnd),
	.combout(\rdata2_M~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~18 .lut_mask = 16'hCEC2;
defparam \rdata2_M~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N12
cycloneive_lcell_comb \rdata2_M~19 (
// Equation(s):
// \rdata2_M~19_combout  = (\rdata2_M[16]~0_combout  & ((\rdata2_M~18_combout  & (\wdat_WB[8]~45_combout )) # (!\rdata2_M~18_combout  & ((ramiframload_8))))) # (!\rdata2_M[16]~0_combout  & (((\rdata2_M~18_combout ))))

	.dataa(\wdat_WB[8]~45_combout ),
	.datab(\dpif.dmemload [8]),
	.datac(\rdata2_M[16]~0_combout ),
	.datad(\rdata2_M~18_combout ),
	.cin(gnd),
	.combout(\rdata2_M~19_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~19 .lut_mask = 16'hAFC0;
defparam \rdata2_M~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N14
cycloneive_lcell_comb \pc_plus_4_EX~8 (
// Equation(s):
// \pc_plus_4_EX~8_combout  = (pc_plus_4_D[9] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[9]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~8_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~8 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N15
dffeas \pc_plus_4_EX[9] (
	.clk(CLK),
	.d(\pc_plus_4_EX~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[9]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[9] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N22
cycloneive_lcell_comb \pc_plus_4_M~8 (
// Equation(s):
// \pc_plus_4_M~8_combout  = (pc_plus_4_EX[9] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_plus_4_EX[9]),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~8_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~8 .lut_mask = 16'h00F0;
defparam \pc_plus_4_M~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N23
dffeas \pc_plus_4_M[9] (
	.clk(CLK),
	.d(\pc_plus_4_M~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[9]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[9] .is_wysiwyg = "true";
defparam \pc_plus_4_M[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N29
dffeas \pc_plus_4_WB[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[9]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[9]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[9] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N12
cycloneive_lcell_comb \dmemload_WB[9]~feeder (
// Equation(s):
// \dmemload_WB[9]~feeder_combout  = ramiframload_9

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(\dmemload_WB[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \dmemload_WB[9]~feeder .lut_mask = 16'hFF00;
defparam \dmemload_WB[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N13
dffeas \dmemload_WB[9] (
	.clk(CLK),
	.d(\dmemload_WB[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[9]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[9] .is_wysiwyg = "true";
defparam \dmemload_WB[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N11
dffeas \porto_WB[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_9),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[9]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[9] .is_wysiwyg = "true";
defparam \porto_WB[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N10
cycloneive_lcell_comb \wdat_WB[9]~42 (
// Equation(s):
// \wdat_WB[9]~42_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[9])) # (!\memToReg_WB~q  & ((porto_WB[9])))))

	.dataa(\jal_WB~q ),
	.datab(dmemload_WB[9]),
	.datac(porto_WB[9]),
	.datad(\memToReg_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[9]~42_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[9]~42 .lut_mask = 16'h4450;
defparam \wdat_WB[9]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N28
cycloneive_lcell_comb \wdat_WB[9]~43 (
// Equation(s):
// \wdat_WB[9]~43_combout  = (!\lui_WB~q  & ((\wdat_WB[9]~42_combout ) # ((\jal_WB~q  & pc_plus_4_WB[9]))))

	.dataa(\jal_WB~q ),
	.datab(\lui_WB~q ),
	.datac(pc_plus_4_WB[9]),
	.datad(\wdat_WB[9]~42_combout ),
	.cin(gnd),
	.combout(\wdat_WB[9]~43_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[9]~43 .lut_mask = 16'h3320;
defparam \wdat_WB[9]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N8
cycloneive_lcell_comb \sw_forwarding_output~20 (
// Equation(s):
// \sw_forwarding_output~20_combout  = (!\lui_M~q  & porto_M_9)

	.dataa(\lui_M~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(porto_M_9),
	.cin(gnd),
	.combout(\sw_forwarding_output~20_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~20 .lut_mask = 16'h5500;
defparam \sw_forwarding_output~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N2
cycloneive_lcell_comb \instruction_D~90 (
// Equation(s):
// \instruction_D~90_combout  = (\branch_or_jump~1_combout  & (ramiframload_9 & iwait))

	.dataa(\branch_or_jump~1_combout ),
	.datab(ramiframload_9),
	.datac(iwait),
	.datad(gnd),
	.cin(gnd),
	.combout(\instruction_D~90_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~90 .lut_mask = 16'h8080;
defparam \instruction_D~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N3
dffeas \instruction_D[9] (
	.clk(CLK),
	.d(\instruction_D~90_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[9]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[9] .is_wysiwyg = "true";
defparam \instruction_D[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N16
cycloneive_lcell_comb \imm_EX~4 (
// Equation(s):
// \imm_EX~4_combout  = (instruction_D[9] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(instruction_D[9]),
	.datac(\branch_taken~0_combout ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\imm_EX~4_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~4 .lut_mask = 16'h8400;
defparam \imm_EX~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N17
dffeas \imm_EX[9] (
	.clk(CLK),
	.d(\imm_EX~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[9]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[9] .is_wysiwyg = "true";
defparam \imm_EX[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N6
cycloneive_lcell_comb \portB~71 (
// Equation(s):
// \portB~71_combout  = (\Equal3~2_combout  & (((\wdat_WB[9]~43_combout ) # (\portB~14_combout )))) # (!\Equal3~2_combout  & (rdata2_EX[9] & ((!\portB~14_combout ))))

	.dataa(rdata2_EX[9]),
	.datab(\wdat_WB[9]~43_combout ),
	.datac(\Equal3~2_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~71_combout ),
	.cout());
// synopsys translate_off
defparam \portB~71 .lut_mask = 16'hF0CA;
defparam \portB~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N2
cycloneive_lcell_comb \portB~72 (
// Equation(s):
// \portB~72_combout  = (\portB~14_combout  & ((\portB~71_combout  & (\sw_forwarding_output~20_combout )) # (!\portB~71_combout  & ((imm_EX[9]))))) # (!\portB~14_combout  & (((\portB~71_combout ))))

	.dataa(\sw_forwarding_output~20_combout ),
	.datab(imm_EX[9]),
	.datac(\portB~14_combout ),
	.datad(\portB~71_combout ),
	.cin(gnd),
	.combout(\portB~72_combout ),
	.cout());
// synopsys translate_off
defparam \portB~72 .lut_mask = 16'hAFC0;
defparam \portB~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N20
cycloneive_lcell_comb \portB~73 (
// Equation(s):
// \portB~73_combout  = (\portB~72_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\ShiftOp_EX~q ),
	.datad(\portB~72_combout ),
	.cin(gnd),
	.combout(\portB~73_combout ),
	.cout());
// synopsys translate_off
defparam \portB~73 .lut_mask = 16'hAF00;
defparam \portB~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N2
cycloneive_lcell_comb \rdata2_EX~40 (
// Equation(s):
// \rdata2_EX~40_combout  = (instruction_D[20] & ((Mux54))) # (!instruction_D[20] & (Mux541))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux54~19_combout ),
	.datad(\REGISTER_FILE|Mux54~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~40_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~40 .lut_mask = 16'hFC30;
defparam \rdata2_EX~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N16
cycloneive_lcell_comb \rdata2_EX~41 (
// Equation(s):
// \rdata2_EX~41_combout  = (\always2~2_combout  & ((\rdata2_EX~40_combout ))) # (!\always2~2_combout  & (\portB~73_combout ))

	.dataa(gnd),
	.datab(\portB~73_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~40_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~41_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~41 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N17
dffeas \rdata2_EX[9] (
	.clk(CLK),
	.d(\rdata2_EX~41_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[9]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[9] .is_wysiwyg = "true";
defparam \rdata2_EX[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N30
cycloneive_lcell_comb \rdata2_M~20 (
// Equation(s):
// \rdata2_M~20_combout  = (\rdata2_M[16]~1_combout  & (\rdata2_M[16]~0_combout )) # (!\rdata2_M[16]~1_combout  & ((\rdata2_M[16]~0_combout  & ((ramiframload_9))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[9]))))

	.dataa(\rdata2_M[16]~1_combout ),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(rdata2_EX[9]),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(\rdata2_M~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~20 .lut_mask = 16'hDC98;
defparam \rdata2_M~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N20
cycloneive_lcell_comb \rdata2_M~21 (
// Equation(s):
// \rdata2_M~21_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~20_combout  & (\wdat_WB[9]~43_combout )) # (!\rdata2_M~20_combout  & ((\sw_forwarding_output~20_combout ))))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~20_combout ))))

	.dataa(\wdat_WB[9]~43_combout ),
	.datab(\sw_forwarding_output~20_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\rdata2_M~20_combout ),
	.cin(gnd),
	.combout(\rdata2_M~21_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~21 .lut_mask = 16'hAFC0;
defparam \rdata2_M~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N18
cycloneive_lcell_comb \pc_plus_4_EX~11 (
// Equation(s):
// \pc_plus_4_EX~11_combout  = (pc_plus_4_D[10] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[10]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~11_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~11 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N19
dffeas \pc_plus_4_EX[10] (
	.clk(CLK),
	.d(\pc_plus_4_EX~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[10]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[10] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N22
cycloneive_lcell_comb \pc_plus_4_M~11 (
// Equation(s):
// \pc_plus_4_M~11_combout  = (pc_plus_4_EX[10] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[10]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~11_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~11 .lut_mask = 16'h00CC;
defparam \pc_plus_4_M~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N23
dffeas \pc_plus_4_M[10] (
	.clk(CLK),
	.d(\pc_plus_4_M~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[10]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[10] .is_wysiwyg = "true";
defparam \pc_plus_4_M[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N3
dffeas \pc_plus_4_WB[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[10]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[10]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[10] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N21
dffeas \porto_WB[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_10),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[10]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[10] .is_wysiwyg = "true";
defparam \porto_WB[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N20
cycloneive_lcell_comb \wdat_WB[10]~48 (
// Equation(s):
// \wdat_WB[10]~48_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[10])) # (!\memToReg_WB~q  & ((porto_WB[10])))))

	.dataa(dmemload_WB[10]),
	.datab(\jal_WB~q ),
	.datac(porto_WB[10]),
	.datad(\memToReg_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[10]~48_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[10]~48 .lut_mask = 16'h2230;
defparam \wdat_WB[10]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N2
cycloneive_lcell_comb \wdat_WB[10]~49 (
// Equation(s):
// \wdat_WB[10]~49_combout  = (!\lui_WB~q  & ((\wdat_WB[10]~48_combout ) # ((\jal_WB~q  & pc_plus_4_WB[10]))))

	.dataa(\lui_WB~q ),
	.datab(\jal_WB~q ),
	.datac(pc_plus_4_WB[10]),
	.datad(\wdat_WB[10]~48_combout ),
	.cin(gnd),
	.combout(\wdat_WB[10]~49_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[10]~49 .lut_mask = 16'h5540;
defparam \wdat_WB[10]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N8
cycloneive_lcell_comb \sw_forwarding_output~23 (
// Equation(s):
// \sw_forwarding_output~23_combout  = (porto_M_10 & !\lui_M~q )

	.dataa(gnd),
	.datab(porto_M_10),
	.datac(gnd),
	.datad(\lui_M~q ),
	.cin(gnd),
	.combout(\sw_forwarding_output~23_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~23 .lut_mask = 16'h00CC;
defparam \sw_forwarding_output~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N18
cycloneive_lcell_comb \rdata2_M~22 (
// Equation(s):
// \rdata2_M~22_combout  = (\rdata2_M[16]~1_combout  & (((\sw_forwarding_output~23_combout ) # (\rdata2_M[16]~0_combout )))) # (!\rdata2_M[16]~1_combout  & (rdata2_EX[10] & ((!\rdata2_M[16]~0_combout ))))

	.dataa(rdata2_EX[10]),
	.datab(\sw_forwarding_output~23_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\rdata2_M[16]~0_combout ),
	.cin(gnd),
	.combout(\rdata2_M~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~22 .lut_mask = 16'hF0CA;
defparam \rdata2_M~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N2
cycloneive_lcell_comb \rdata2_M~23 (
// Equation(s):
// \rdata2_M~23_combout  = (\rdata2_M~22_combout  & ((\wdat_WB[10]~49_combout ) # ((!\rdata2_M[16]~0_combout )))) # (!\rdata2_M~22_combout  & (((ramiframload_10 & \rdata2_M[16]~0_combout ))))

	.dataa(\wdat_WB[10]~49_combout ),
	.datab(\rdata2_M~22_combout ),
	.datac(\dpif.dmemload [10]),
	.datad(\rdata2_M[16]~0_combout ),
	.cin(gnd),
	.combout(\rdata2_M~23_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~23 .lut_mask = 16'hB8CC;
defparam \rdata2_M~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N16
cycloneive_lcell_comb \sw_forwarding_output~22 (
// Equation(s):
// \sw_forwarding_output~22_combout  = (!\lui_M~q  & porto_M_11)

	.dataa(gnd),
	.datab(gnd),
	.datac(\lui_M~q ),
	.datad(porto_M_11),
	.cin(gnd),
	.combout(\sw_forwarding_output~22_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~22 .lut_mask = 16'h0F00;
defparam \sw_forwarding_output~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N4
cycloneive_lcell_comb \pc_plus_4_EX~10 (
// Equation(s):
// \pc_plus_4_EX~10_combout  = (pc_plus_4_D[11] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(pc_plus_4_D[11]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\branch_taken~0_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~10_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~10 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N5
dffeas \pc_plus_4_EX[11] (
	.clk(CLK),
	.d(\pc_plus_4_EX~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[11]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[11] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N20
cycloneive_lcell_comb \pc_plus_4_M~10 (
// Equation(s):
// \pc_plus_4_M~10_combout  = (pc_plus_4_EX[11] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[11]),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_plus_4_M~10_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~10 .lut_mask = 16'h0C0C;
defparam \pc_plus_4_M~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N21
dffeas \pc_plus_4_M[11] (
	.clk(CLK),
	.d(\pc_plus_4_M~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[11]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[11] .is_wysiwyg = "true";
defparam \pc_plus_4_M[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N19
dffeas \pc_plus_4_WB[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[11]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[11]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[11] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N21
dffeas \porto_WB[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_11),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[11]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[11] .is_wysiwyg = "true";
defparam \porto_WB[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N20
cycloneive_lcell_comb \wdat_WB[11]~46 (
// Equation(s):
// \wdat_WB[11]~46_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[11])) # (!\memToReg_WB~q  & ((porto_WB[11])))))

	.dataa(dmemload_WB[11]),
	.datab(\memToReg_WB~q ),
	.datac(porto_WB[11]),
	.datad(\jal_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[11]~46_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[11]~46 .lut_mask = 16'h00B8;
defparam \wdat_WB[11]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N18
cycloneive_lcell_comb \wdat_WB[11]~47 (
// Equation(s):
// \wdat_WB[11]~47_combout  = (!\lui_WB~q  & ((\wdat_WB[11]~46_combout ) # ((\jal_WB~q  & pc_plus_4_WB[11]))))

	.dataa(\jal_WB~q ),
	.datab(\lui_WB~q ),
	.datac(pc_plus_4_WB[11]),
	.datad(\wdat_WB[11]~46_combout ),
	.cin(gnd),
	.combout(\wdat_WB[11]~47_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[11]~47 .lut_mask = 16'h3320;
defparam \wdat_WB[11]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N20
cycloneive_lcell_comb \rdata2_M~24 (
// Equation(s):
// \rdata2_M~24_combout  = (\rdata2_M[16]~0_combout  & (((ramiframload_11) # (\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[11] & ((!\rdata2_M[16]~1_combout ))))

	.dataa(rdata2_EX[11]),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\dpif.dmemload [11]),
	.datad(\rdata2_M[16]~1_combout ),
	.cin(gnd),
	.combout(\rdata2_M~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~24 .lut_mask = 16'hCCE2;
defparam \rdata2_M~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N6
cycloneive_lcell_comb \rdata2_M~25 (
// Equation(s):
// \rdata2_M~25_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~24_combout  & ((\wdat_WB[11]~47_combout ))) # (!\rdata2_M~24_combout  & (\sw_forwarding_output~22_combout )))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~24_combout ))))

	.dataa(\sw_forwarding_output~22_combout ),
	.datab(\rdata2_M[16]~1_combout ),
	.datac(\wdat_WB[11]~47_combout ),
	.datad(\rdata2_M~24_combout ),
	.cin(gnd),
	.combout(\rdata2_M~25_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~25 .lut_mask = 16'hF388;
defparam \rdata2_M~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N6
cycloneive_lcell_comb \rdata2_EX~38 (
// Equation(s):
// \rdata2_EX~38_combout  = (instruction_D[20] & ((Mux51))) # (!instruction_D[20] & (Mux511))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux51~19_combout ),
	.datad(\REGISTER_FILE|Mux51~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~38_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~38 .lut_mask = 16'hFA50;
defparam \rdata2_EX~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N2
cycloneive_lcell_comb \rdata2_EX~39 (
// Equation(s):
// \rdata2_EX~39_combout  = (\always2~2_combout  & ((\rdata2_EX~38_combout ))) # (!\always2~2_combout  & (\portB~70_combout ))

	.dataa(\portB~70_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~38_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~39_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~39 .lut_mask = 16'hFA0A;
defparam \rdata2_EX~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N3
dffeas \rdata2_EX[12] (
	.clk(CLK),
	.d(\rdata2_EX~39_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[12]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[12] .is_wysiwyg = "true";
defparam \rdata2_EX[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N24
cycloneive_lcell_comb \sw_forwarding_output~19 (
// Equation(s):
// \sw_forwarding_output~19_combout  = (!\lui_M~q  & porto_M_12)

	.dataa(\lui_M~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(porto_M_12),
	.cin(gnd),
	.combout(\sw_forwarding_output~19_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~19 .lut_mask = 16'h5500;
defparam \sw_forwarding_output~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N22
cycloneive_lcell_comb \rdata2_M~26 (
// Equation(s):
// \rdata2_M~26_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & ((\rdata2_M[16]~1_combout  & ((\sw_forwarding_output~19_combout ))) # (!\rdata2_M[16]~1_combout  & (rdata2_EX[12]))))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(rdata2_EX[12]),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\sw_forwarding_output~19_combout ),
	.cin(gnd),
	.combout(\rdata2_M~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~26 .lut_mask = 16'hF4A4;
defparam \rdata2_M~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N17
dffeas \dmemload_WB[12] (
	.clk(CLK),
	.d(\dpif.dmemload [12]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[12]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[12] .is_wysiwyg = "true";
defparam \dmemload_WB[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N19
dffeas \porto_WB[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_12),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[12]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[12] .is_wysiwyg = "true";
defparam \porto_WB[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N18
cycloneive_lcell_comb \wdat_WB[12]~40 (
// Equation(s):
// \wdat_WB[12]~40_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[12])) # (!\memToReg_WB~q  & ((porto_WB[12])))))

	.dataa(\memToReg_WB~q ),
	.datab(dmemload_WB[12]),
	.datac(porto_WB[12]),
	.datad(\jal_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[12]~40_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[12]~40 .lut_mask = 16'h00D8;
defparam \wdat_WB[12]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N8
cycloneive_lcell_comb \pc_plus_4_M~13 (
// Equation(s):
// \pc_plus_4_M~13_combout  = (pc_plus_4_EX[12] & !\wsel_M~0_combout )

	.dataa(pc_plus_4_EX[12]),
	.datab(gnd),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~13_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~13 .lut_mask = 16'h00AA;
defparam \pc_plus_4_M~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N9
dffeas \pc_plus_4_M[12] (
	.clk(CLK),
	.d(\pc_plus_4_M~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[12]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[12] .is_wysiwyg = "true";
defparam \pc_plus_4_M[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N21
dffeas \pc_plus_4_WB[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[12]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[12]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[12] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N20
cycloneive_lcell_comb \wdat_WB[12]~41 (
// Equation(s):
// \wdat_WB[12]~41_combout  = (!\lui_WB~q  & ((\wdat_WB[12]~40_combout ) # ((\jal_WB~q  & pc_plus_4_WB[12]))))

	.dataa(\jal_WB~q ),
	.datab(\wdat_WB[12]~40_combout ),
	.datac(pc_plus_4_WB[12]),
	.datad(\lui_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[12]~41_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[12]~41 .lut_mask = 16'h00EC;
defparam \wdat_WB[12]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N22
cycloneive_lcell_comb \rdata2_M~27 (
// Equation(s):
// \rdata2_M~27_combout  = (\rdata2_M~26_combout  & ((\wdat_WB[12]~41_combout ) # ((!\rdata2_M[16]~0_combout )))) # (!\rdata2_M~26_combout  & (((\rdata2_M[16]~0_combout  & ramiframload_12))))

	.dataa(\rdata2_M~26_combout ),
	.datab(\wdat_WB[12]~41_combout ),
	.datac(\rdata2_M[16]~0_combout ),
	.datad(\dpif.dmemload [12]),
	.cin(gnd),
	.combout(\rdata2_M~27_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~27 .lut_mask = 16'hDA8A;
defparam \rdata2_M~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N30
cycloneive_lcell_comb \sw_forwarding_output~18 (
// Equation(s):
// \sw_forwarding_output~18_combout  = (porto_M_13 & !\lui_M~q )

	.dataa(gnd),
	.datab(gnd),
	.datac(porto_M_13),
	.datad(\lui_M~q ),
	.cin(gnd),
	.combout(\sw_forwarding_output~18_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~18 .lut_mask = 16'h00F0;
defparam \sw_forwarding_output~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N16
cycloneive_lcell_comb \pc_plus_4_EX~12 (
// Equation(s):
// \pc_plus_4_EX~12_combout  = (pc_plus_4_D[13] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[13]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~12_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~12 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y36_N17
dffeas \pc_plus_4_EX[13] (
	.clk(CLK),
	.d(\pc_plus_4_EX~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[13]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[13] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N22
cycloneive_lcell_comb \pc_plus_4_M~12 (
// Equation(s):
// \pc_plus_4_M~12_combout  = (pc_plus_4_EX[13] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_plus_4_EX[13]),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~12_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~12 .lut_mask = 16'h00F0;
defparam \pc_plus_4_M~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N23
dffeas \pc_plus_4_M[13] (
	.clk(CLK),
	.d(\pc_plus_4_M~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[13]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[13] .is_wysiwyg = "true";
defparam \pc_plus_4_M[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N29
dffeas \pc_plus_4_WB[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[13]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[13]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[13] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N3
dffeas \dmemload_WB[13] (
	.clk(CLK),
	.d(\dpif.dmemload [13]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[13]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[13] .is_wysiwyg = "true";
defparam \dmemload_WB[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N7
dffeas \porto_WB[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_13),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[13]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[13] .is_wysiwyg = "true";
defparam \porto_WB[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N6
cycloneive_lcell_comb \wdat_WB[13]~38 (
// Equation(s):
// \wdat_WB[13]~38_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[13])) # (!\memToReg_WB~q  & ((porto_WB[13])))))

	.dataa(\memToReg_WB~q ),
	.datab(dmemload_WB[13]),
	.datac(porto_WB[13]),
	.datad(\jal_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[13]~38_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[13]~38 .lut_mask = 16'h00D8;
defparam \wdat_WB[13]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N28
cycloneive_lcell_comb \wdat_WB[13]~39 (
// Equation(s):
// \wdat_WB[13]~39_combout  = (!\lui_WB~q  & ((\wdat_WB[13]~38_combout ) # ((\jal_WB~q  & pc_plus_4_WB[13]))))

	.dataa(\jal_WB~q ),
	.datab(\lui_WB~q ),
	.datac(pc_plus_4_WB[13]),
	.datad(\wdat_WB[13]~38_combout ),
	.cin(gnd),
	.combout(\wdat_WB[13]~39_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[13]~39 .lut_mask = 16'h3320;
defparam \wdat_WB[13]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N20
cycloneive_lcell_comb \rdata2_M~28 (
// Equation(s):
// \rdata2_M~28_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout ) # (ramiframload_13)))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[13] & (!\rdata2_M[16]~1_combout )))

	.dataa(rdata2_EX[13]),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\dpif.dmemload [13]),
	.cin(gnd),
	.combout(\rdata2_M~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~28 .lut_mask = 16'hCEC2;
defparam \rdata2_M~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N8
cycloneive_lcell_comb \rdata2_M~29 (
// Equation(s):
// \rdata2_M~29_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~28_combout  & ((\wdat_WB[13]~39_combout ))) # (!\rdata2_M~28_combout  & (\sw_forwarding_output~18_combout )))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~28_combout ))))

	.dataa(\sw_forwarding_output~18_combout ),
	.datab(\wdat_WB[13]~39_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\rdata2_M~28_combout ),
	.cin(gnd),
	.combout(\rdata2_M~29_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~29 .lut_mask = 16'hCFA0;
defparam \rdata2_M~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N16
cycloneive_lcell_comb \instruction_D~87 (
// Equation(s):
// \instruction_D~87_combout  = (iwait & (\branch_or_jump~1_combout  & ramiframload_14))

	.dataa(iwait),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\dpif.dmemload [14]),
	.cin(gnd),
	.combout(\instruction_D~87_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~87 .lut_mask = 16'hA000;
defparam \instruction_D~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N17
dffeas \instruction_D[14] (
	.clk(CLK),
	.d(\instruction_D~87_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[14]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[14] .is_wysiwyg = "true";
defparam \instruction_D[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N26
cycloneive_lcell_comb \imm_EX~1 (
// Equation(s):
// \imm_EX~1_combout  = (\branch_or_jump~2_combout  & (instruction_D[14] & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(instruction_D[14]),
	.datac(\branch_taken~0_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\imm_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~1 .lut_mask = 16'h8008;
defparam \imm_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N27
dffeas \imm_EX[14] (
	.clk(CLK),
	.d(\imm_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[14]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[14] .is_wysiwyg = "true";
defparam \imm_EX[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N4
cycloneive_lcell_comb \portB~65 (
// Equation(s):
// \portB~65_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & (imm_EX[14])) # (!\portB~14_combout  & ((rdata2_EX[14])))))

	.dataa(\ShiftOp_EX~q ),
	.datab(imm_EX[14]),
	.datac(rdata2_EX[14]),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~65_combout ),
	.cout());
// synopsys translate_off
defparam \portB~65 .lut_mask = 16'h4450;
defparam \portB~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N2
cycloneive_lcell_comb \portB~111 (
// Equation(s):
// \portB~111_combout  = (\portB~14_combout  & (((!\lui_M~q  & porto_M_14)))) # (!\portB~14_combout  & (\wdat_WB[14]~37_combout ))

	.dataa(\wdat_WB[14]~37_combout ),
	.datab(\lui_M~q ),
	.datac(porto_M_14),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~111_combout ),
	.cout());
// synopsys translate_off
defparam \portB~111 .lut_mask = 16'h30AA;
defparam \portB~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N30
cycloneive_lcell_comb \portB~66 (
// Equation(s):
// \portB~66_combout  = (\Equal3~2_combout  & ((\portB~111_combout ))) # (!\Equal3~2_combout  & (\portB~65_combout ))

	.dataa(\Equal3~2_combout ),
	.datab(\portB~65_combout ),
	.datac(gnd),
	.datad(\portB~111_combout ),
	.cin(gnd),
	.combout(\portB~66_combout ),
	.cout());
// synopsys translate_off
defparam \portB~66 .lut_mask = 16'hEE44;
defparam \portB~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N10
cycloneive_lcell_comb \rdata2_EX~34 (
// Equation(s):
// \rdata2_EX~34_combout  = (instruction_D[20] & (Mux49)) # (!instruction_D[20] & ((Mux491)))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux49~9_combout ),
	.datad(\REGISTER_FILE|Mux49~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~34_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~34 .lut_mask = 16'hF3C0;
defparam \rdata2_EX~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N26
cycloneive_lcell_comb \rdata2_EX~35 (
// Equation(s):
// \rdata2_EX~35_combout  = (\always2~2_combout  & ((\rdata2_EX~34_combout ))) # (!\always2~2_combout  & (\portB~66_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portB~66_combout ),
	.datad(\rdata2_EX~34_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~35_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~35 .lut_mask = 16'hFC30;
defparam \rdata2_EX~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N27
dffeas \rdata2_EX[14] (
	.clk(CLK),
	.d(\rdata2_EX~35_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[14]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[14] .is_wysiwyg = "true";
defparam \rdata2_EX[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N6
cycloneive_lcell_comb \rdata2_M~30 (
// Equation(s):
// \rdata2_M~30_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & ((\rdata2_M[16]~1_combout  & (\sw_forwarding_output~17_combout )) # (!\rdata2_M[16]~1_combout  & ((rdata2_EX[14])))))

	.dataa(\sw_forwarding_output~17_combout ),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(rdata2_EX[14]),
	.cin(gnd),
	.combout(\rdata2_M~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~30 .lut_mask = 16'hE3E0;
defparam \rdata2_M~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N20
cycloneive_lcell_comb \pc_plus_4_M~15 (
// Equation(s):
// \pc_plus_4_M~15_combout  = (pc_plus_4_EX[14] & !\wsel_M~0_combout )

	.dataa(pc_plus_4_EX[14]),
	.datab(gnd),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~15_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~15 .lut_mask = 16'h00AA;
defparam \pc_plus_4_M~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N21
dffeas \pc_plus_4_M[14] (
	.clk(CLK),
	.d(\pc_plus_4_M~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[14]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[14] .is_wysiwyg = "true";
defparam \pc_plus_4_M[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N13
dffeas \pc_plus_4_WB[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[14]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[14]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[14] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N7
dffeas \porto_WB[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_14),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[14]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[14] .is_wysiwyg = "true";
defparam \porto_WB[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N6
cycloneive_lcell_comb \wdat_WB[14]~36 (
// Equation(s):
// \wdat_WB[14]~36_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[14])) # (!\memToReg_WB~q  & ((porto_WB[14])))))

	.dataa(dmemload_WB[14]),
	.datab(\memToReg_WB~q ),
	.datac(porto_WB[14]),
	.datad(\jal_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[14]~36_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[14]~36 .lut_mask = 16'h00B8;
defparam \wdat_WB[14]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N12
cycloneive_lcell_comb \wdat_WB[14]~37 (
// Equation(s):
// \wdat_WB[14]~37_combout  = (!\lui_WB~q  & ((\wdat_WB[14]~36_combout ) # ((\jal_WB~q  & pc_plus_4_WB[14]))))

	.dataa(\jal_WB~q ),
	.datab(\lui_WB~q ),
	.datac(pc_plus_4_WB[14]),
	.datad(\wdat_WB[14]~36_combout ),
	.cin(gnd),
	.combout(\wdat_WB[14]~37_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[14]~37 .lut_mask = 16'h3320;
defparam \wdat_WB[14]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N24
cycloneive_lcell_comb \rdata2_M~31 (
// Equation(s):
// \rdata2_M~31_combout  = (\rdata2_M~30_combout  & ((\wdat_WB[14]~37_combout ) # ((!\rdata2_M[16]~0_combout )))) # (!\rdata2_M~30_combout  & (((\rdata2_M[16]~0_combout  & ramiframload_14))))

	.dataa(\rdata2_M~30_combout ),
	.datab(\wdat_WB[14]~37_combout ),
	.datac(\rdata2_M[16]~0_combout ),
	.datad(\dpif.dmemload [14]),
	.cin(gnd),
	.combout(\rdata2_M~31_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~31 .lut_mask = 16'hDA8A;
defparam \rdata2_M~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N16
cycloneive_lcell_comb \pc_plus_4_M~14 (
// Equation(s):
// \pc_plus_4_M~14_combout  = (pc_plus_4_EX[15] & !\wsel_M~0_combout )

	.dataa(pc_plus_4_EX[15]),
	.datab(gnd),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~14_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~14 .lut_mask = 16'h00AA;
defparam \pc_plus_4_M~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N17
dffeas \pc_plus_4_M[15] (
	.clk(CLK),
	.d(\pc_plus_4_M~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[15]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[15] .is_wysiwyg = "true";
defparam \pc_plus_4_M[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N17
dffeas \pc_plus_4_WB[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[15]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[15]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[15] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N3
dffeas \porto_WB[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_15),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[15]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[15] .is_wysiwyg = "true";
defparam \porto_WB[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N2
cycloneive_lcell_comb \wdat_WB[15]~34 (
// Equation(s):
// \wdat_WB[15]~34_combout  = (!\jal_WB~q  & ((\memToReg_WB~q  & (dmemload_WB[15])) # (!\memToReg_WB~q  & ((porto_WB[15])))))

	.dataa(dmemload_WB[15]),
	.datab(\jal_WB~q ),
	.datac(porto_WB[15]),
	.datad(\memToReg_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[15]~34_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[15]~34 .lut_mask = 16'h2230;
defparam \wdat_WB[15]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N16
cycloneive_lcell_comb \wdat_WB[15]~35 (
// Equation(s):
// \wdat_WB[15]~35_combout  = (!\lui_WB~q  & ((\wdat_WB[15]~34_combout ) # ((\jal_WB~q  & pc_plus_4_WB[15]))))

	.dataa(\jal_WB~q ),
	.datab(\lui_WB~q ),
	.datac(pc_plus_4_WB[15]),
	.datad(\wdat_WB[15]~34_combout ),
	.cin(gnd),
	.combout(\wdat_WB[15]~35_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[15]~35 .lut_mask = 16'h3320;
defparam \wdat_WB[15]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N2
cycloneive_lcell_comb \instruction_D~86 (
// Equation(s):
// \instruction_D~86_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_15))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(iwait),
	.datad(ramiframload_15),
	.cin(gnd),
	.combout(\instruction_D~86_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~86 .lut_mask = 16'hA000;
defparam \instruction_D~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N3
dffeas \instruction_D[15] (
	.clk(CLK),
	.d(\instruction_D~86_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[15]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[15] .is_wysiwyg = "true";
defparam \instruction_D[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N30
cycloneive_lcell_comb \imm_EX~0 (
// Equation(s):
// \imm_EX~0_combout  = (instruction_D[15] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_taken~0_combout ),
	.datab(instruction_D[15]),
	.datac(\branch_or_jump~2_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\imm_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~0 .lut_mask = 16'h8040;
defparam \imm_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N31
dffeas \imm_EX[15] (
	.clk(CLK),
	.d(\imm_EX~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[15]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[15] .is_wysiwyg = "true";
defparam \imm_EX[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N22
cycloneive_lcell_comb \portB~63 (
// Equation(s):
// \portB~63_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & ((imm_EX[15]))) # (!\portB~14_combout  & (rdata2_EX[15]))))

	.dataa(rdata2_EX[15]),
	.datab(\ShiftOp_EX~q ),
	.datac(imm_EX[15]),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~63_combout ),
	.cout());
// synopsys translate_off
defparam \portB~63 .lut_mask = 16'h3022;
defparam \portB~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N10
cycloneive_lcell_comb \portB~110 (
// Equation(s):
// \portB~110_combout  = (\portB~14_combout  & (porto_M_15 & ((!\lui_M~q )))) # (!\portB~14_combout  & (((\wdat_WB[15]~35_combout ))))

	.dataa(porto_M_15),
	.datab(\wdat_WB[15]~35_combout ),
	.datac(\lui_M~q ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~110_combout ),
	.cout());
// synopsys translate_off
defparam \portB~110 .lut_mask = 16'h0ACC;
defparam \portB~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N14
cycloneive_lcell_comb \portB~64 (
// Equation(s):
// \portB~64_combout  = (\Equal3~2_combout  & ((\portB~110_combout ))) # (!\Equal3~2_combout  & (\portB~63_combout ))

	.dataa(gnd),
	.datab(\Equal3~2_combout ),
	.datac(\portB~63_combout ),
	.datad(\portB~110_combout ),
	.cin(gnd),
	.combout(\portB~64_combout ),
	.cout());
// synopsys translate_off
defparam \portB~64 .lut_mask = 16'hFC30;
defparam \portB~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N28
cycloneive_lcell_comb \rdata2_EX~32 (
// Equation(s):
// \rdata2_EX~32_combout  = (instruction_D[20] & (Mux48)) # (!instruction_D[20] & ((Mux481)))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux48~9_combout ),
	.datad(\REGISTER_FILE|Mux48~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~32_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~32 .lut_mask = 16'hF3C0;
defparam \rdata2_EX~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N8
cycloneive_lcell_comb \rdata2_EX~33 (
// Equation(s):
// \rdata2_EX~33_combout  = (\always2~2_combout  & ((\rdata2_EX~32_combout ))) # (!\always2~2_combout  & (\portB~64_combout ))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\portB~64_combout ),
	.datad(\rdata2_EX~32_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~33_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~33 .lut_mask = 16'hFC30;
defparam \rdata2_EX~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y29_N9
dffeas \rdata2_EX[15] (
	.clk(CLK),
	.d(\rdata2_EX~33_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[15]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[15] .is_wysiwyg = "true";
defparam \rdata2_EX[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N4
cycloneive_lcell_comb \rdata2_M~32 (
// Equation(s):
// \rdata2_M~32_combout  = (\rdata2_M[16]~1_combout  & (((\rdata2_M[16]~0_combout )))) # (!\rdata2_M[16]~1_combout  & ((\rdata2_M[16]~0_combout  & (ramiframload_15)) # (!\rdata2_M[16]~0_combout  & ((rdata2_EX[15])))))

	.dataa(\rdata2_M[16]~1_combout ),
	.datab(ramiframload_15),
	.datac(\rdata2_M[16]~0_combout ),
	.datad(rdata2_EX[15]),
	.cin(gnd),
	.combout(\rdata2_M~32_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~32 .lut_mask = 16'hE5E0;
defparam \rdata2_M~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N16
cycloneive_lcell_comb \sw_forwarding_output~16 (
// Equation(s):
// \sw_forwarding_output~16_combout  = (!\lui_M~q  & porto_M_15)

	.dataa(gnd),
	.datab(gnd),
	.datac(\lui_M~q ),
	.datad(porto_M_15),
	.cin(gnd),
	.combout(\sw_forwarding_output~16_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~16 .lut_mask = 16'h0F00;
defparam \sw_forwarding_output~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N20
cycloneive_lcell_comb \rdata2_M~33 (
// Equation(s):
// \rdata2_M~33_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~32_combout  & (\wdat_WB[15]~35_combout )) # (!\rdata2_M~32_combout  & ((\sw_forwarding_output~16_combout ))))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~32_combout ))))

	.dataa(\wdat_WB[15]~35_combout ),
	.datab(\rdata2_M[16]~1_combout ),
	.datac(\rdata2_M~32_combout ),
	.datad(\sw_forwarding_output~16_combout ),
	.cin(gnd),
	.combout(\rdata2_M~33_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~33 .lut_mask = 16'hBCB0;
defparam \rdata2_M~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N17
dffeas \dmemload_WB[16] (
	.clk(CLK),
	.d(\dpif.dmemload [16]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[16]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[16] .is_wysiwyg = "true";
defparam \dmemload_WB[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N30
cycloneive_lcell_comb \instruction_D~81 (
// Equation(s):
// \instruction_D~81_combout  = (\branch_or_jump~1_combout  & (ramiframload_0 & iwait))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(\dpif.dmemload [0]),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~81_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~81 .lut_mask = 16'hA000;
defparam \instruction_D~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N31
dffeas \instruction_D[0] (
	.clk(CLK),
	.d(\instruction_D~81_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[0]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[0] .is_wysiwyg = "true";
defparam \instruction_D[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N18
cycloneive_lcell_comb \imm_EX~11 (
// Equation(s):
// \imm_EX~11_combout  = (\branch_or_jump~2_combout  & (instruction_D[0] & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(\branch_taken~0_combout ),
	.datac(instruction_D[0]),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\imm_EX~11_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~11 .lut_mask = 16'h8020;
defparam \imm_EX~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N1
dffeas \imm_EX[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\imm_EX~11_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[0]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[0] .is_wysiwyg = "true";
defparam \imm_EX[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N22
cycloneive_lcell_comb \imm_M~15 (
// Equation(s):
// \imm_M~15_combout  = (!\wsel_M~0_combout  & imm_EX[0])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(imm_EX[0]),
	.cin(gnd),
	.combout(\imm_M~15_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~15 .lut_mask = 16'h0F00;
defparam \imm_M~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N23
dffeas \imm_M[0] (
	.clk(CLK),
	.d(\imm_M~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[0]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[0] .is_wysiwyg = "true";
defparam \imm_M[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N19
dffeas \imm_WB[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[0]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[0]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[0] .is_wysiwyg = "true";
defparam \imm_WB[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N12
cycloneive_lcell_comb \wdat_WB[28]~1 (
// Equation(s):
// \wdat_WB[28]~1_combout  = (\lui_WB~q ) # ((!\jal_WB~q  & \memToReg_WB~q ))

	.dataa(\jal_WB~q ),
	.datab(\memToReg_WB~q ),
	.datac(gnd),
	.datad(\lui_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[28]~1_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[28]~1 .lut_mask = 16'hFF44;
defparam \wdat_WB[28]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N29
dffeas \porto_WB[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_16),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[16]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[16] .is_wysiwyg = "true";
defparam \porto_WB[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N8
cycloneive_lcell_comb \wdat_WB[28]~0 (
// Equation(s):
// \wdat_WB[28]~0_combout  = (\jal_WB~q ) # (\lui_WB~q )

	.dataa(\jal_WB~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\lui_WB~q ),
	.cin(gnd),
	.combout(\wdat_WB[28]~0_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[28]~0 .lut_mask = 16'hFFAA;
defparam \wdat_WB[28]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N28
cycloneive_lcell_comb \wdat_WB[16]~32 (
// Equation(s):
// \wdat_WB[16]~32_combout  = (\wdat_WB[28]~1_combout  & (((\wdat_WB[28]~0_combout )))) # (!\wdat_WB[28]~1_combout  & ((\wdat_WB[28]~0_combout  & (pc_plus_4_WB[16])) # (!\wdat_WB[28]~0_combout  & ((porto_WB[16])))))

	.dataa(pc_plus_4_WB[16]),
	.datab(\wdat_WB[28]~1_combout ),
	.datac(porto_WB[16]),
	.datad(\wdat_WB[28]~0_combout ),
	.cin(gnd),
	.combout(\wdat_WB[16]~32_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[16]~32 .lut_mask = 16'hEE30;
defparam \wdat_WB[16]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N18
cycloneive_lcell_comb \wdat_WB[16]~33 (
// Equation(s):
// \wdat_WB[16]~33_combout  = (\wdat_WB[28]~1_combout  & ((\wdat_WB[16]~32_combout  & ((imm_WB[0]))) # (!\wdat_WB[16]~32_combout  & (dmemload_WB[16])))) # (!\wdat_WB[28]~1_combout  & (((\wdat_WB[16]~32_combout ))))

	.dataa(\wdat_WB[28]~1_combout ),
	.datab(dmemload_WB[16]),
	.datac(imm_WB[0]),
	.datad(\wdat_WB[16]~32_combout ),
	.cin(gnd),
	.combout(\wdat_WB[16]~33_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[16]~33 .lut_mask = 16'hF588;
defparam \wdat_WB[16]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N20
cycloneive_lcell_comb \sw_forwarding_output~15 (
// Equation(s):
// \sw_forwarding_output~15_combout  = (\lui_M~q  & ((imm_M[0]))) # (!\lui_M~q  & (porto_M_16))

	.dataa(gnd),
	.datab(\lui_M~q ),
	.datac(porto_M_16),
	.datad(imm_M[0]),
	.cin(gnd),
	.combout(\sw_forwarding_output~15_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~15 .lut_mask = 16'hFC30;
defparam \sw_forwarding_output~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N22
cycloneive_lcell_comb \rdata2_EX~30 (
// Equation(s):
// \rdata2_EX~30_combout  = (instruction_D[20] & (Mux47)) # (!instruction_D[20] & ((Mux471)))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux47~9_combout ),
	.datad(\REGISTER_FILE|Mux47~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~30 .lut_mask = 16'hF3C0;
defparam \rdata2_EX~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N2
cycloneive_lcell_comb \portB~61 (
// Equation(s):
// \portB~61_combout  = (\portB~14_combout  & (\sw_forwarding_output~15_combout )) # (!\portB~14_combout  & ((\wdat_WB[16]~33_combout )))

	.dataa(gnd),
	.datab(\sw_forwarding_output~15_combout ),
	.datac(\portB~14_combout ),
	.datad(\wdat_WB[16]~33_combout ),
	.cin(gnd),
	.combout(\portB~61_combout ),
	.cout());
// synopsys translate_off
defparam \portB~61 .lut_mask = 16'hCFC0;
defparam \portB~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N22
cycloneive_lcell_comb \portB~62 (
// Equation(s):
// \portB~62_combout  = (\Equal3~2_combout  & ((\portB~61_combout ))) # (!\Equal3~2_combout  & (\portB~60_combout ))

	.dataa(\portB~60_combout ),
	.datab(\Equal3~2_combout ),
	.datac(gnd),
	.datad(\portB~61_combout ),
	.cin(gnd),
	.combout(\portB~62_combout ),
	.cout());
// synopsys translate_off
defparam \portB~62 .lut_mask = 16'hEE22;
defparam \portB~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N24
cycloneive_lcell_comb \rdata2_EX~31 (
// Equation(s):
// \rdata2_EX~31_combout  = (\always2~2_combout  & (\rdata2_EX~30_combout )) # (!\always2~2_combout  & ((\portB~62_combout )))

	.dataa(gnd),
	.datab(\always2~2_combout ),
	.datac(\rdata2_EX~30_combout ),
	.datad(\portB~62_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~31_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~31 .lut_mask = 16'hF3C0;
defparam \rdata2_EX~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N25
dffeas \rdata2_EX[16] (
	.clk(CLK),
	.d(\rdata2_EX~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[16]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[16] .is_wysiwyg = "true";
defparam \rdata2_EX[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N26
cycloneive_lcell_comb \rdata2_M~34 (
// Equation(s):
// \rdata2_M~34_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & ((\rdata2_M[16]~1_combout  & (\sw_forwarding_output~15_combout )) # (!\rdata2_M[16]~1_combout  & ((rdata2_EX[16])))))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(\sw_forwarding_output~15_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(rdata2_EX[16]),
	.cin(gnd),
	.combout(\rdata2_M~34_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~34 .lut_mask = 16'hE5E0;
defparam \rdata2_M~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N10
cycloneive_lcell_comb \rdata2_M~35 (
// Equation(s):
// \rdata2_M~35_combout  = (\rdata2_M[16]~0_combout  & ((\rdata2_M~34_combout  & ((\wdat_WB[16]~33_combout ))) # (!\rdata2_M~34_combout  & (ramiframload_16)))) # (!\rdata2_M[16]~0_combout  & (((\rdata2_M~34_combout ))))

	.dataa(\dpif.dmemload [16]),
	.datab(\wdat_WB[16]~33_combout ),
	.datac(\rdata2_M[16]~0_combout ),
	.datad(\rdata2_M~34_combout ),
	.cin(gnd),
	.combout(\rdata2_M~35_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~35 .lut_mask = 16'hCFA0;
defparam \rdata2_M~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N0
cycloneive_lcell_comb \pc_plus_4[17]~30 (
// Equation(s):
// \pc_plus_4[17]~30_combout  = (pc_out_17 & (!\pc_plus_4[16]~29 )) # (!pc_out_17 & ((\pc_plus_4[16]~29 ) # (GND)))
// \pc_plus_4[17]~31  = CARRY((!\pc_plus_4[16]~29 ) # (!pc_out_17))

	.dataa(pc_out_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[16]~29 ),
	.combout(\pc_plus_4[17]~30_combout ),
	.cout(\pc_plus_4[17]~31 ));
// synopsys translate_off
defparam \pc_plus_4[17]~30 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[17]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N20
cycloneive_lcell_comb \pc_plus_4_D~16 (
// Equation(s):
// \pc_plus_4_D~16_combout  = (\pc_plus_4[17]~30_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(iwait),
	.datab(gnd),
	.datac(\pc_plus_4[17]~30_combout ),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~16_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~16 .lut_mask = 16'hA0F0;
defparam \pc_plus_4_D~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N21
dffeas \pc_plus_4_D[17] (
	.clk(CLK),
	.d(\pc_plus_4_D~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[17]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[17] .is_wysiwyg = "true";
defparam \pc_plus_4_D[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N14
cycloneive_lcell_comb \pc_plus_4_EX~16 (
// Equation(s):
// \pc_plus_4_EX~16_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[17] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_D[17]),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~16_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~16 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N15
dffeas \pc_plus_4_EX[17] (
	.clk(CLK),
	.d(\pc_plus_4_EX~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[17]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[17] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N14
cycloneive_lcell_comb \pc_plus_4_M~16 (
// Equation(s):
// \pc_plus_4_M~16_combout  = (!\wsel_M~0_combout  & pc_plus_4_EX[17])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(pc_plus_4_EX[17]),
	.cin(gnd),
	.combout(\pc_plus_4_M~16_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~16 .lut_mask = 16'h0F00;
defparam \pc_plus_4_M~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N15
dffeas \pc_plus_4_M[17] (
	.clk(CLK),
	.d(\pc_plus_4_M~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[17]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[17] .is_wysiwyg = "true";
defparam \pc_plus_4_M[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N13
dffeas \pc_plus_4_WB[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[17]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[17]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[17] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N3
dffeas \porto_WB[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_17),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[17]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[17] .is_wysiwyg = "true";
defparam \porto_WB[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N2
cycloneive_lcell_comb \wdat_WB[17]~30 (
// Equation(s):
// \wdat_WB[17]~30_combout  = (\wdat_WB[28]~0_combout  & (((\wdat_WB[28]~1_combout )))) # (!\wdat_WB[28]~0_combout  & ((\wdat_WB[28]~1_combout  & (dmemload_WB[17])) # (!\wdat_WB[28]~1_combout  & ((porto_WB[17])))))

	.dataa(dmemload_WB[17]),
	.datab(\wdat_WB[28]~0_combout ),
	.datac(porto_WB[17]),
	.datad(\wdat_WB[28]~1_combout ),
	.cin(gnd),
	.combout(\wdat_WB[17]~30_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[17]~30 .lut_mask = 16'hEE30;
defparam \wdat_WB[17]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N12
cycloneive_lcell_comb \wdat_WB[17]~31 (
// Equation(s):
// \wdat_WB[17]~31_combout  = (\wdat_WB[28]~0_combout  & ((\wdat_WB[17]~30_combout  & (imm_WB[1])) # (!\wdat_WB[17]~30_combout  & ((pc_plus_4_WB[17]))))) # (!\wdat_WB[28]~0_combout  & (((\wdat_WB[17]~30_combout ))))

	.dataa(imm_WB[1]),
	.datab(\wdat_WB[28]~0_combout ),
	.datac(pc_plus_4_WB[17]),
	.datad(\wdat_WB[17]~30_combout ),
	.cin(gnd),
	.combout(\wdat_WB[17]~31_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[17]~31 .lut_mask = 16'hBBC0;
defparam \wdat_WB[17]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N30
cycloneive_lcell_comb \instruction_D~84 (
// Equation(s):
// \instruction_D~84_combout  = (\branch_or_jump~1_combout  & (ramiframload_1 & iwait))

	.dataa(\branch_or_jump~1_combout ),
	.datab(\dpif.dmemload [1]),
	.datac(iwait),
	.datad(gnd),
	.cin(gnd),
	.combout(\instruction_D~84_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~84 .lut_mask = 16'h8080;
defparam \instruction_D~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N31
dffeas \instruction_D[1] (
	.clk(CLK),
	.d(\instruction_D~84_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[1]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[1] .is_wysiwyg = "true";
defparam \instruction_D[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N14
cycloneive_lcell_comb \imm_EX~12 (
// Equation(s):
// \imm_EX~12_combout  = (instruction_D[1] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(\branch_taken~0_combout ),
	.datac(instruction_D[1]),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\imm_EX~12_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~12 .lut_mask = 16'h9000;
defparam \imm_EX~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N15
dffeas \imm_EX[1] (
	.clk(CLK),
	.d(\imm_EX~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[1]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[1] .is_wysiwyg = "true";
defparam \imm_EX[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N14
cycloneive_lcell_comb \imm_M~14 (
// Equation(s):
// \imm_M~14_combout  = (!\wsel_M~0_combout  & imm_EX[1])

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(imm_EX[1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\imm_M~14_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~14 .lut_mask = 16'h3030;
defparam \imm_M~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y32_N15
dffeas \imm_M[1] (
	.clk(CLK),
	.d(\imm_M~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[1]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[1] .is_wysiwyg = "true";
defparam \imm_M[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N26
cycloneive_lcell_comb \sw_forwarding_output~14 (
// Equation(s):
// \sw_forwarding_output~14_combout  = (\lui_M~q  & (imm_M[1])) # (!\lui_M~q  & ((porto_M_17)))

	.dataa(\lui_M~q ),
	.datab(gnd),
	.datac(imm_M[1]),
	.datad(porto_M_17),
	.cin(gnd),
	.combout(\sw_forwarding_output~14_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~14 .lut_mask = 16'hF5A0;
defparam \sw_forwarding_output~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N20
cycloneive_lcell_comb \rdata2_EX~28 (
// Equation(s):
// \rdata2_EX~28_combout  = (instruction_D[20] & ((Mux46))) # (!instruction_D[20] & (Mux461))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux46~19_combout ),
	.datad(\REGISTER_FILE|Mux46~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~28 .lut_mask = 16'hFC30;
defparam \rdata2_EX~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N14
cycloneive_lcell_comb \rdata2_EX~29 (
// Equation(s):
// \rdata2_EX~29_combout  = (\always2~2_combout  & ((\rdata2_EX~28_combout ))) # (!\always2~2_combout  & (\portB~59_combout ))

	.dataa(\portB~59_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~28_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~29_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~29 .lut_mask = 16'hFA0A;
defparam \rdata2_EX~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N15
dffeas \rdata2_EX[17] (
	.clk(CLK),
	.d(\rdata2_EX~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[17]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[17] .is_wysiwyg = "true";
defparam \rdata2_EX[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N10
cycloneive_lcell_comb \rdata2_M~36 (
// Equation(s):
// \rdata2_M~36_combout  = (\rdata2_M[16]~0_combout  & ((ramiframload_17) # ((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & (((rdata2_EX[17] & !\rdata2_M[16]~1_combout ))))

	.dataa(\dpif.dmemload [17]),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(rdata2_EX[17]),
	.datad(\rdata2_M[16]~1_combout ),
	.cin(gnd),
	.combout(\rdata2_M~36_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~36 .lut_mask = 16'hCCB8;
defparam \rdata2_M~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N24
cycloneive_lcell_comb \rdata2_M~37 (
// Equation(s):
// \rdata2_M~37_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~36_combout  & (\wdat_WB[17]~31_combout )) # (!\rdata2_M~36_combout  & ((\sw_forwarding_output~14_combout ))))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~36_combout ))))

	.dataa(\wdat_WB[17]~31_combout ),
	.datab(\rdata2_M[16]~1_combout ),
	.datac(\sw_forwarding_output~14_combout ),
	.datad(\rdata2_M~36_combout ),
	.cin(gnd),
	.combout(\rdata2_M~37_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~37 .lut_mask = 16'hBBC0;
defparam \rdata2_M~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N22
cycloneive_lcell_comb \imm_EX~13 (
// Equation(s):
// \imm_EX~13_combout  = (\branch_or_jump~2_combout  & (instruction_D[2] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(\branch_or_jump~2_combout ),
	.datac(\branch_taken~0_combout ),
	.datad(instruction_D[2]),
	.cin(gnd),
	.combout(\imm_EX~13_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~13 .lut_mask = 16'h8400;
defparam \imm_EX~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N23
dffeas \imm_EX[2] (
	.clk(CLK),
	.d(\imm_EX~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[2]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[2] .is_wysiwyg = "true";
defparam \imm_EX[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N6
cycloneive_lcell_comb \imm_M~13 (
// Equation(s):
// \imm_M~13_combout  = (imm_EX[2] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(imm_EX[2]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\imm_M~13_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~13 .lut_mask = 16'h00CC;
defparam \imm_M~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y35_N7
dffeas \imm_M[2] (
	.clk(CLK),
	.d(\imm_M~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[2]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[2] .is_wysiwyg = "true";
defparam \imm_M[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N17
dffeas \imm_WB[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[2]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[2]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[2] .is_wysiwyg = "true";
defparam \imm_WB[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N3
dffeas \porto_WB[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_18),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[18]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[18] .is_wysiwyg = "true";
defparam \porto_WB[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N2
cycloneive_lcell_comb \wdat_WB[18]~28 (
// Equation(s):
// \wdat_WB[18]~28_combout  = (\wdat_WB[28]~1_combout  & (((\wdat_WB[28]~0_combout )))) # (!\wdat_WB[28]~1_combout  & ((\wdat_WB[28]~0_combout  & (pc_plus_4_WB[18])) # (!\wdat_WB[28]~0_combout  & ((porto_WB[18])))))

	.dataa(pc_plus_4_WB[18]),
	.datab(\wdat_WB[28]~1_combout ),
	.datac(porto_WB[18]),
	.datad(\wdat_WB[28]~0_combout ),
	.cin(gnd),
	.combout(\wdat_WB[18]~28_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[18]~28 .lut_mask = 16'hEE30;
defparam \wdat_WB[18]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N16
cycloneive_lcell_comb \wdat_WB[18]~29 (
// Equation(s):
// \wdat_WB[18]~29_combout  = (\wdat_WB[28]~1_combout  & ((\wdat_WB[18]~28_combout  & ((imm_WB[2]))) # (!\wdat_WB[18]~28_combout  & (dmemload_WB[18])))) # (!\wdat_WB[28]~1_combout  & (((\wdat_WB[18]~28_combout ))))

	.dataa(dmemload_WB[18]),
	.datab(\wdat_WB[28]~1_combout ),
	.datac(imm_WB[2]),
	.datad(\wdat_WB[18]~28_combout ),
	.cin(gnd),
	.combout(\wdat_WB[18]~29_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[18]~29 .lut_mask = 16'hF388;
defparam \wdat_WB[18]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N12
cycloneive_lcell_comb \sw_forwarding_output~13 (
// Equation(s):
// \sw_forwarding_output~13_combout  = (\lui_M~q  & (imm_M[2])) # (!\lui_M~q  & ((porto_M_18)))

	.dataa(imm_M[2]),
	.datab(porto_M_18),
	.datac(\lui_M~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\sw_forwarding_output~13_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~13 .lut_mask = 16'hACAC;
defparam \sw_forwarding_output~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N22
cycloneive_lcell_comb \portB~55 (
// Equation(s):
// \portB~55_combout  = (\portB~14_combout  & ((\sw_forwarding_output~13_combout ))) # (!\portB~14_combout  & (\wdat_WB[18]~29_combout ))

	.dataa(gnd),
	.datab(\wdat_WB[18]~29_combout ),
	.datac(\sw_forwarding_output~13_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~55_combout ),
	.cout());
// synopsys translate_off
defparam \portB~55 .lut_mask = 16'hF0CC;
defparam \portB~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N0
cycloneive_lcell_comb \portB~54 (
// Equation(s):
// \portB~54_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & (\sign_ext[16]~0_combout )) # (!\portB~14_combout  & ((rdata2_EX[18])))))

	.dataa(\sign_ext[16]~0_combout ),
	.datab(rdata2_EX[18]),
	.datac(\ShiftOp_EX~q ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~54_combout ),
	.cout());
// synopsys translate_off
defparam \portB~54 .lut_mask = 16'h0A0C;
defparam \portB~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N24
cycloneive_lcell_comb \portB~56 (
// Equation(s):
// \portB~56_combout  = (\Equal3~2_combout  & (\portB~55_combout )) # (!\Equal3~2_combout  & ((\portB~54_combout )))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~55_combout ),
	.datad(\portB~54_combout ),
	.cin(gnd),
	.combout(\portB~56_combout ),
	.cout());
// synopsys translate_off
defparam \portB~56 .lut_mask = 16'hF5A0;
defparam \portB~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N28
cycloneive_lcell_comb \rdata2_EX~26 (
// Equation(s):
// \rdata2_EX~26_combout  = (instruction_D[20] & ((Mux45))) # (!instruction_D[20] & (Mux451))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux45~19_combout ),
	.datad(\REGISTER_FILE|Mux45~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~26 .lut_mask = 16'hFC30;
defparam \rdata2_EX~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N0
cycloneive_lcell_comb \rdata2_EX~27 (
// Equation(s):
// \rdata2_EX~27_combout  = (\always2~2_combout  & ((\rdata2_EX~26_combout ))) # (!\always2~2_combout  & (\portB~56_combout ))

	.dataa(gnd),
	.datab(\portB~56_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~26_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~27_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~27 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N1
dffeas \rdata2_EX[18] (
	.clk(CLK),
	.d(\rdata2_EX~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[18]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[18] .is_wysiwyg = "true";
defparam \rdata2_EX[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N4
cycloneive_lcell_comb \rdata2_M~38 (
// Equation(s):
// \rdata2_M~38_combout  = (\rdata2_M[16]~1_combout  & (((\sw_forwarding_output~13_combout ) # (\rdata2_M[16]~0_combout )))) # (!\rdata2_M[16]~1_combout  & (rdata2_EX[18] & ((!\rdata2_M[16]~0_combout ))))

	.dataa(\rdata2_M[16]~1_combout ),
	.datab(rdata2_EX[18]),
	.datac(\sw_forwarding_output~13_combout ),
	.datad(\rdata2_M[16]~0_combout ),
	.cin(gnd),
	.combout(\rdata2_M~38_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~38 .lut_mask = 16'hAAE4;
defparam \rdata2_M~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N16
cycloneive_lcell_comb \rdata2_M~39 (
// Equation(s):
// \rdata2_M~39_combout  = (\rdata2_M[16]~0_combout  & ((\rdata2_M~38_combout  & (\wdat_WB[18]~29_combout )) # (!\rdata2_M~38_combout  & ((ramiframload_18))))) # (!\rdata2_M[16]~0_combout  & (((\rdata2_M~38_combout ))))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(\wdat_WB[18]~29_combout ),
	.datac(\rdata2_M~38_combout ),
	.datad(ramiframload_18),
	.cin(gnd),
	.combout(\rdata2_M~39_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~39 .lut_mask = 16'hDAD0;
defparam \rdata2_M~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N8
cycloneive_lcell_comb \imm_EX~14 (
// Equation(s):
// \imm_EX~14_combout  = (\branch_or_jump~2_combout  & (instruction_D[3] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(\branch_or_jump~2_combout ),
	.datac(instruction_D[3]),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\imm_EX~14_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~14 .lut_mask = 16'h8040;
defparam \imm_EX~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N9
dffeas \imm_EX[3] (
	.clk(CLK),
	.d(\imm_EX~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[3]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[3] .is_wysiwyg = "true";
defparam \imm_EX[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N8
cycloneive_lcell_comb \imm_M~12 (
// Equation(s):
// \imm_M~12_combout  = (imm_EX[3] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(imm_EX[3]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\imm_M~12_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~12 .lut_mask = 16'h00CC;
defparam \imm_M~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N9
dffeas \imm_M[3] (
	.clk(CLK),
	.d(\imm_M~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[3]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[3] .is_wysiwyg = "true";
defparam \imm_M[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N14
cycloneive_lcell_comb \sw_forwarding_output~12 (
// Equation(s):
// \sw_forwarding_output~12_combout  = (\lui_M~q  & (imm_M[3])) # (!\lui_M~q  & ((porto_M_19)))

	.dataa(gnd),
	.datab(imm_M[3]),
	.datac(porto_M_19),
	.datad(\lui_M~q ),
	.cin(gnd),
	.combout(\sw_forwarding_output~12_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~12 .lut_mask = 16'hCCF0;
defparam \sw_forwarding_output~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N14
cycloneive_lcell_comb \imm_WB[3]~feeder (
// Equation(s):
// \imm_WB[3]~feeder_combout  = imm_M[3]

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(imm_M[3]),
	.cin(gnd),
	.combout(\imm_WB[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \imm_WB[3]~feeder .lut_mask = 16'hFF00;
defparam \imm_WB[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N15
dffeas \imm_WB[3] (
	.clk(CLK),
	.d(\imm_WB[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[3]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[3] .is_wysiwyg = "true";
defparam \imm_WB[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N4
cycloneive_lcell_comb \pc_plus_4[19]~34 (
// Equation(s):
// \pc_plus_4[19]~34_combout  = (pc_out_19 & (!\pc_plus_4[18]~33 )) # (!pc_out_19 & ((\pc_plus_4[18]~33 ) # (GND)))
// \pc_plus_4[19]~35  = CARRY((!\pc_plus_4[18]~33 ) # (!pc_out_19))

	.dataa(pc_out_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[18]~33 ),
	.combout(\pc_plus_4[19]~34_combout ),
	.cout(\pc_plus_4[19]~35 ));
// synopsys translate_off
defparam \pc_plus_4[19]~34 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[19]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N26
cycloneive_lcell_comb \pc_plus_4_D~18 (
// Equation(s):
// \pc_plus_4_D~18_combout  = (\pc_plus_4[19]~34_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(\pc_plus_4[19]~34_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~18_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~18 .lut_mask = 16'hF300;
defparam \pc_plus_4_D~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N27
dffeas \pc_plus_4_D[19] (
	.clk(CLK),
	.d(\pc_plus_4_D~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[19]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[19] .is_wysiwyg = "true";
defparam \pc_plus_4_D[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N2
cycloneive_lcell_comb \pc_plus_4_EX~18 (
// Equation(s):
// \pc_plus_4_EX~18_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[19] & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(\branch_taken~0_combout ),
	.datac(pc_plus_4_D[19]),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~18_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~18 .lut_mask = 16'h8020;
defparam \pc_plus_4_EX~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N3
dffeas \pc_plus_4_EX[19] (
	.clk(CLK),
	.d(\pc_plus_4_EX~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[19]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[19] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N18
cycloneive_lcell_comb \pc_plus_4_M~18 (
// Equation(s):
// \pc_plus_4_M~18_combout  = (!\wsel_M~0_combout  & pc_plus_4_EX[19])

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(gnd),
	.datad(pc_plus_4_EX[19]),
	.cin(gnd),
	.combout(\pc_plus_4_M~18_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~18 .lut_mask = 16'h3300;
defparam \pc_plus_4_M~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N19
dffeas \pc_plus_4_M[19] (
	.clk(CLK),
	.d(\pc_plus_4_M~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[19]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[19] .is_wysiwyg = "true";
defparam \pc_plus_4_M[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N5
dffeas \pc_plus_4_WB[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[19]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[19]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[19] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N1
dffeas \porto_WB[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_19),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[19]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[19] .is_wysiwyg = "true";
defparam \porto_WB[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N0
cycloneive_lcell_comb \wdat_WB[19]~26 (
// Equation(s):
// \wdat_WB[19]~26_combout  = (\wdat_WB[28]~1_combout  & ((dmemload_WB[19]) # ((\wdat_WB[28]~0_combout )))) # (!\wdat_WB[28]~1_combout  & (((porto_WB[19] & !\wdat_WB[28]~0_combout ))))

	.dataa(dmemload_WB[19]),
	.datab(\wdat_WB[28]~1_combout ),
	.datac(porto_WB[19]),
	.datad(\wdat_WB[28]~0_combout ),
	.cin(gnd),
	.combout(\wdat_WB[19]~26_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[19]~26 .lut_mask = 16'hCCB8;
defparam \wdat_WB[19]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N4
cycloneive_lcell_comb \wdat_WB[19]~27 (
// Equation(s):
// \wdat_WB[19]~27_combout  = (\wdat_WB[28]~0_combout  & ((\wdat_WB[19]~26_combout  & (imm_WB[3])) # (!\wdat_WB[19]~26_combout  & ((pc_plus_4_WB[19]))))) # (!\wdat_WB[28]~0_combout  & (((\wdat_WB[19]~26_combout ))))

	.dataa(\wdat_WB[28]~0_combout ),
	.datab(imm_WB[3]),
	.datac(pc_plus_4_WB[19]),
	.datad(\wdat_WB[19]~26_combout ),
	.cin(gnd),
	.combout(\wdat_WB[19]~27_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[19]~27 .lut_mask = 16'hDDA0;
defparam \wdat_WB[19]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N26
cycloneive_lcell_comb \portB~51 (
// Equation(s):
// \portB~51_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & (\sign_ext[16]~0_combout )) # (!\portB~14_combout  & ((rdata2_EX[19])))))

	.dataa(\sign_ext[16]~0_combout ),
	.datab(\ShiftOp_EX~q ),
	.datac(rdata2_EX[19]),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~51_combout ),
	.cout());
// synopsys translate_off
defparam \portB~51 .lut_mask = 16'h2230;
defparam \portB~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N28
cycloneive_lcell_comb \portB~52 (
// Equation(s):
// \portB~52_combout  = (\portB~14_combout  & (\sw_forwarding_output~12_combout )) # (!\portB~14_combout  & ((\wdat_WB[19]~27_combout )))

	.dataa(gnd),
	.datab(\sw_forwarding_output~12_combout ),
	.datac(\wdat_WB[19]~27_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~52_combout ),
	.cout());
// synopsys translate_off
defparam \portB~52 .lut_mask = 16'hCCF0;
defparam \portB~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N14
cycloneive_lcell_comb \portB~53 (
// Equation(s):
// \portB~53_combout  = (\Equal3~2_combout  & ((\portB~52_combout ))) # (!\Equal3~2_combout  & (\portB~51_combout ))

	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(\portB~51_combout ),
	.datad(\portB~52_combout ),
	.cin(gnd),
	.combout(\portB~53_combout ),
	.cout());
// synopsys translate_off
defparam \portB~53 .lut_mask = 16'hFA50;
defparam \portB~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N6
cycloneive_lcell_comb \rdata2_EX~24 (
// Equation(s):
// \rdata2_EX~24_combout  = (instruction_D[20] & (Mux44)) # (!instruction_D[20] & ((Mux441)))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux44~9_combout ),
	.datad(\REGISTER_FILE|Mux44~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~24 .lut_mask = 16'hF3C0;
defparam \rdata2_EX~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N18
cycloneive_lcell_comb \rdata2_EX~25 (
// Equation(s):
// \rdata2_EX~25_combout  = (\always2~2_combout  & ((\rdata2_EX~24_combout ))) # (!\always2~2_combout  & (\portB~53_combout ))

	.dataa(gnd),
	.datab(\portB~53_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~24_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~25_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~25 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N19
dffeas \rdata2_EX[19] (
	.clk(CLK),
	.d(\rdata2_EX~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[19]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[19] .is_wysiwyg = "true";
defparam \rdata2_EX[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N16
cycloneive_lcell_comb \rdata2_M~40 (
// Equation(s):
// \rdata2_M~40_combout  = (\rdata2_M[16]~0_combout  & ((ramiframload_19) # ((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & (((rdata2_EX[19] & !\rdata2_M[16]~1_combout ))))

	.dataa(ramiframload_19),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(rdata2_EX[19]),
	.datad(\rdata2_M[16]~1_combout ),
	.cin(gnd),
	.combout(\rdata2_M~40_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~40 .lut_mask = 16'hCCB8;
defparam \rdata2_M~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N2
cycloneive_lcell_comb \rdata2_M~41 (
// Equation(s):
// \rdata2_M~41_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~40_combout  & ((\wdat_WB[19]~27_combout ))) # (!\rdata2_M~40_combout  & (\sw_forwarding_output~12_combout )))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~40_combout ))))

	.dataa(\sw_forwarding_output~12_combout ),
	.datab(\rdata2_M[16]~1_combout ),
	.datac(\wdat_WB[19]~27_combout ),
	.datad(\rdata2_M~40_combout ),
	.cin(gnd),
	.combout(\rdata2_M~41_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~41 .lut_mask = 16'hF388;
defparam \rdata2_M~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N28
cycloneive_lcell_comb \sw_forwarding_output~11 (
// Equation(s):
// \sw_forwarding_output~11_combout  = (\lui_M~q  & (imm_M[4])) # (!\lui_M~q  & ((porto_M_20)))

	.dataa(imm_M[4]),
	.datab(porto_M_20),
	.datac(gnd),
	.datad(\lui_M~q ),
	.cin(gnd),
	.combout(\sw_forwarding_output~11_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~11 .lut_mask = 16'hAACC;
defparam \sw_forwarding_output~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N4
cycloneive_lcell_comb \rdata2_M~42 (
// Equation(s):
// \rdata2_M~42_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & ((\rdata2_M[16]~1_combout  & ((\sw_forwarding_output~11_combout ))) # (!\rdata2_M[16]~1_combout  & (rdata2_EX[20]))))

	.dataa(rdata2_EX[20]),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\sw_forwarding_output~11_combout ),
	.cin(gnd),
	.combout(\rdata2_M~42_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~42 .lut_mask = 16'hF2C2;
defparam \rdata2_M~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N29
dffeas \dmemload_WB[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_20),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[20]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[20] .is_wysiwyg = "true";
defparam \dmemload_WB[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N12
cycloneive_lcell_comb \imm_M~11 (
// Equation(s):
// \imm_M~11_combout  = (!\wsel_M~0_combout  & imm_EX[4])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(imm_EX[4]),
	.cin(gnd),
	.combout(\imm_M~11_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~11 .lut_mask = 16'h0F00;
defparam \imm_M~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N13
dffeas \imm_M[4] (
	.clk(CLK),
	.d(\imm_M~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[4]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[4] .is_wysiwyg = "true";
defparam \imm_M[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N11
dffeas \imm_WB[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[4]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[4]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[4] .is_wysiwyg = "true";
defparam \imm_WB[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N6
cycloneive_lcell_comb \pc_plus_4[20]~36 (
// Equation(s):
// \pc_plus_4[20]~36_combout  = (pc_out_20 & (\pc_plus_4[19]~35  $ (GND))) # (!pc_out_20 & (!\pc_plus_4[19]~35  & VCC))
// \pc_plus_4[20]~37  = CARRY((pc_out_20 & !\pc_plus_4[19]~35 ))

	.dataa(gnd),
	.datab(pc_out_20),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[19]~35 ),
	.combout(\pc_plus_4[20]~36_combout ),
	.cout(\pc_plus_4[20]~37 ));
// synopsys translate_off
defparam \pc_plus_4[20]~36 .lut_mask = 16'hC30C;
defparam \pc_plus_4[20]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N4
cycloneive_lcell_comb \pc_plus_4_D~21 (
// Equation(s):
// \pc_plus_4_D~21_combout  = (\pc_plus_4[20]~36_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(iwait),
	.datab(\branch_or_jump~1_combout ),
	.datac(gnd),
	.datad(\pc_plus_4[20]~36_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~21_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~21 .lut_mask = 16'hBB00;
defparam \pc_plus_4_D~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N5
dffeas \pc_plus_4_D[20] (
	.clk(CLK),
	.d(\pc_plus_4_D~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[20]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[20] .is_wysiwyg = "true";
defparam \pc_plus_4_D[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N14
cycloneive_lcell_comb \pc_plus_4_EX~21 (
// Equation(s):
// \pc_plus_4_EX~21_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[20] & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_D[20]),
	.datac(\branch_taken~0_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~21_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~21 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N15
dffeas \pc_plus_4_EX[20] (
	.clk(CLK),
	.d(\pc_plus_4_EX~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[20]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[20] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N8
cycloneive_lcell_comb \pc_plus_4_M~21 (
// Equation(s):
// \pc_plus_4_M~21_combout  = (pc_plus_4_EX[20] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[20]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~21_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~21 .lut_mask = 16'h00CC;
defparam \pc_plus_4_M~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N9
dffeas \pc_plus_4_M[20] (
	.clk(CLK),
	.d(\pc_plus_4_M~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[20]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[20] .is_wysiwyg = "true";
defparam \pc_plus_4_M[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N18
cycloneive_lcell_comb \pc_plus_4_WB[20]~feeder (
// Equation(s):
// \pc_plus_4_WB[20]~feeder_combout  = pc_plus_4_M[20]

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pc_plus_4_M[20]),
	.cin(gnd),
	.combout(\pc_plus_4_WB[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_WB[20]~feeder .lut_mask = 16'hFF00;
defparam \pc_plus_4_WB[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N19
dffeas \pc_plus_4_WB[20] (
	.clk(CLK),
	.d(\pc_plus_4_WB[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[20]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[20] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N21
dffeas \porto_WB[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_20),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[20]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[20] .is_wysiwyg = "true";
defparam \porto_WB[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N20
cycloneive_lcell_comb \wdat_WB[20]~24 (
// Equation(s):
// \wdat_WB[20]~24_combout  = (\wdat_WB[28]~1_combout  & (((\wdat_WB[28]~0_combout )))) # (!\wdat_WB[28]~1_combout  & ((\wdat_WB[28]~0_combout  & (pc_plus_4_WB[20])) # (!\wdat_WB[28]~0_combout  & ((porto_WB[20])))))

	.dataa(\wdat_WB[28]~1_combout ),
	.datab(pc_plus_4_WB[20]),
	.datac(porto_WB[20]),
	.datad(\wdat_WB[28]~0_combout ),
	.cin(gnd),
	.combout(\wdat_WB[20]~24_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[20]~24 .lut_mask = 16'hEE50;
defparam \wdat_WB[20]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N10
cycloneive_lcell_comb \wdat_WB[20]~25 (
// Equation(s):
// \wdat_WB[20]~25_combout  = (\wdat_WB[28]~1_combout  & ((\wdat_WB[20]~24_combout  & ((imm_WB[4]))) # (!\wdat_WB[20]~24_combout  & (dmemload_WB[20])))) # (!\wdat_WB[28]~1_combout  & (((\wdat_WB[20]~24_combout ))))

	.dataa(\wdat_WB[28]~1_combout ),
	.datab(dmemload_WB[20]),
	.datac(imm_WB[4]),
	.datad(\wdat_WB[20]~24_combout ),
	.cin(gnd),
	.combout(\wdat_WB[20]~25_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[20]~25 .lut_mask = 16'hF588;
defparam \wdat_WB[20]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N0
cycloneive_lcell_comb \rdata2_M~43 (
// Equation(s):
// \rdata2_M~43_combout  = (\rdata2_M~42_combout  & (((\wdat_WB[20]~25_combout ) # (!\rdata2_M[16]~0_combout )))) # (!\rdata2_M~42_combout  & (ramiframload_20 & (\rdata2_M[16]~0_combout )))

	.dataa(ramiframload_20),
	.datab(\rdata2_M~42_combout ),
	.datac(\rdata2_M[16]~0_combout ),
	.datad(\wdat_WB[20]~25_combout ),
	.cin(gnd),
	.combout(\rdata2_M~43_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~43 .lut_mask = 16'hEC2C;
defparam \rdata2_M~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N16
cycloneive_lcell_comb \sw_forwarding_output~10 (
// Equation(s):
// \sw_forwarding_output~10_combout  = (\lui_M~q  & (imm_M[5])) # (!\lui_M~q  & ((porto_M_21)))

	.dataa(imm_M[5]),
	.datab(gnd),
	.datac(\lui_M~q ),
	.datad(porto_M_21),
	.cin(gnd),
	.combout(\sw_forwarding_output~10_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~10 .lut_mask = 16'hAFA0;
defparam \sw_forwarding_output~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N26
cycloneive_lcell_comb \imm_EX~10 (
// Equation(s):
// \imm_EX~10_combout  = (instruction_D[5] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(instruction_D[5]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\branch_taken~0_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\imm_EX~10_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~10 .lut_mask = 16'h8008;
defparam \imm_EX~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N27
dffeas \imm_EX[5] (
	.clk(CLK),
	.d(\imm_EX~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[5]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[5] .is_wysiwyg = "true";
defparam \imm_EX[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N6
cycloneive_lcell_comb \imm_M~10 (
// Equation(s):
// \imm_M~10_combout  = (imm_EX[5] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(imm_EX[5]),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\imm_M~10_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~10 .lut_mask = 16'h0C0C;
defparam \imm_M~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N7
dffeas \imm_M[5] (
	.clk(CLK),
	.d(\imm_M~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[5]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[5] .is_wysiwyg = "true";
defparam \imm_M[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N9
dffeas \imm_WB[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[5]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[5]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[5] .is_wysiwyg = "true";
defparam \imm_WB[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N7
dffeas \porto_WB[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_21),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[21]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[21] .is_wysiwyg = "true";
defparam \porto_WB[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N6
cycloneive_lcell_comb \wdat_WB[21]~22 (
// Equation(s):
// \wdat_WB[21]~22_combout  = (\wdat_WB[28]~0_combout  & (((\wdat_WB[28]~1_combout )))) # (!\wdat_WB[28]~0_combout  & ((\wdat_WB[28]~1_combout  & (dmemload_WB[21])) # (!\wdat_WB[28]~1_combout  & ((porto_WB[21])))))

	.dataa(dmemload_WB[21]),
	.datab(\wdat_WB[28]~0_combout ),
	.datac(porto_WB[21]),
	.datad(\wdat_WB[28]~1_combout ),
	.cin(gnd),
	.combout(\wdat_WB[21]~22_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[21]~22 .lut_mask = 16'hEE30;
defparam \wdat_WB[21]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N14
cycloneive_lcell_comb \wdat_WB[21]~23 (
// Equation(s):
// \wdat_WB[21]~23_combout  = (\wdat_WB[28]~0_combout  & ((\wdat_WB[21]~22_combout  & ((imm_WB[5]))) # (!\wdat_WB[21]~22_combout  & (pc_plus_4_WB[21])))) # (!\wdat_WB[28]~0_combout  & (((\wdat_WB[21]~22_combout ))))

	.dataa(pc_plus_4_WB[21]),
	.datab(imm_WB[5]),
	.datac(\wdat_WB[28]~0_combout ),
	.datad(\wdat_WB[21]~22_combout ),
	.cin(gnd),
	.combout(\wdat_WB[21]~23_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[21]~23 .lut_mask = 16'hCFA0;
defparam \wdat_WB[21]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N30
cycloneive_lcell_comb \ExtOp_EX~1 (
// Equation(s):
// \ExtOp_EX~1_combout  = (\ExtOp_EX~0_combout  & (!instruction_D[28] & WideOr8))

	.dataa(\ExtOp_EX~0_combout ),
	.datab(instruction_D[28]),
	.datac(gnd),
	.datad(\CONTROL_UNIT|WideOr8~0_combout ),
	.cin(gnd),
	.combout(\ExtOp_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \ExtOp_EX~1 .lut_mask = 16'h2200;
defparam \ExtOp_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N31
dffeas ExtOp_EX(
	.clk(CLK),
	.d(\ExtOp_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\ExtOp_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam ExtOp_EX.is_wysiwyg = "true";
defparam ExtOp_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N14
cycloneive_lcell_comb \sign_ext[16]~0 (
// Equation(s):
// \sign_ext[16]~0_combout  = (imm_EX[15] & \ExtOp_EX~q )

	.dataa(gnd),
	.datab(gnd),
	.datac(imm_EX[15]),
	.datad(\ExtOp_EX~q ),
	.cin(gnd),
	.combout(\sign_ext[16]~0_combout ),
	.cout());
// synopsys translate_off
defparam \sign_ext[16]~0 .lut_mask = 16'hF000;
defparam \sign_ext[16]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N22
cycloneive_lcell_comb \portB~45 (
// Equation(s):
// \portB~45_combout  = (!\ShiftOp_EX~q  & ((\portB~14_combout  & ((\sign_ext[16]~0_combout ))) # (!\portB~14_combout  & (rdata2_EX[21]))))

	.dataa(rdata2_EX[21]),
	.datab(\ShiftOp_EX~q ),
	.datac(\sign_ext[16]~0_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~45_combout ),
	.cout());
// synopsys translate_off
defparam \portB~45 .lut_mask = 16'h3022;
defparam \portB~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N24
cycloneive_lcell_comb \portB~46 (
// Equation(s):
// \portB~46_combout  = (\portB~14_combout  & (\sw_forwarding_output~10_combout )) # (!\portB~14_combout  & ((\wdat_WB[21]~23_combout )))

	.dataa(gnd),
	.datab(\sw_forwarding_output~10_combout ),
	.datac(\wdat_WB[21]~23_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~46_combout ),
	.cout());
// synopsys translate_off
defparam \portB~46 .lut_mask = 16'hCCF0;
defparam \portB~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N26
cycloneive_lcell_comb \portB~47 (
// Equation(s):
// \portB~47_combout  = (\Equal3~2_combout  & ((\portB~46_combout ))) # (!\Equal3~2_combout  & (\portB~45_combout ))

	.dataa(gnd),
	.datab(\Equal3~2_combout ),
	.datac(\portB~45_combout ),
	.datad(\portB~46_combout ),
	.cin(gnd),
	.combout(\portB~47_combout ),
	.cout());
// synopsys translate_off
defparam \portB~47 .lut_mask = 16'hFC30;
defparam \portB~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N24
cycloneive_lcell_comb \rdata2_EX~20 (
// Equation(s):
// \rdata2_EX~20_combout  = (instruction_D[20] & ((Mux42))) # (!instruction_D[20] & (Mux421))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux42~19_combout ),
	.datad(\REGISTER_FILE|Mux42~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~20 .lut_mask = 16'hFA50;
defparam \rdata2_EX~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N4
cycloneive_lcell_comb \rdata2_EX~21 (
// Equation(s):
// \rdata2_EX~21_combout  = (\always2~2_combout  & ((\rdata2_EX~20_combout ))) # (!\always2~2_combout  & (\portB~47_combout ))

	.dataa(gnd),
	.datab(\portB~47_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~20_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~21_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~21 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N5
dffeas \rdata2_EX[21] (
	.clk(CLK),
	.d(\rdata2_EX~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[21]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[21] .is_wysiwyg = "true";
defparam \rdata2_EX[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N18
cycloneive_lcell_comb \rdata2_M~44 (
// Equation(s):
// \rdata2_M~44_combout  = (\rdata2_M[16]~1_combout  & (((\rdata2_M[16]~0_combout )))) # (!\rdata2_M[16]~1_combout  & ((\rdata2_M[16]~0_combout  & ((ramiframload_21))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[21]))))

	.dataa(\rdata2_M[16]~1_combout ),
	.datab(rdata2_EX[21]),
	.datac(\dpif.dmemload [21]),
	.datad(\rdata2_M[16]~0_combout ),
	.cin(gnd),
	.combout(\rdata2_M~44_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~44 .lut_mask = 16'hFA44;
defparam \rdata2_M~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N10
cycloneive_lcell_comb \rdata2_M~45 (
// Equation(s):
// \rdata2_M~45_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~44_combout  & ((\wdat_WB[21]~23_combout ))) # (!\rdata2_M~44_combout  & (\sw_forwarding_output~10_combout )))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~44_combout ))))

	.dataa(\rdata2_M[16]~1_combout ),
	.datab(\sw_forwarding_output~10_combout ),
	.datac(\wdat_WB[21]~23_combout ),
	.datad(\rdata2_M~44_combout ),
	.cin(gnd),
	.combout(\rdata2_M~45_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~45 .lut_mask = 16'hF588;
defparam \rdata2_M~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N10
cycloneive_lcell_comb \rdata2_EX~18 (
// Equation(s):
// \rdata2_EX~18_combout  = (instruction_D[20] & ((Mux41))) # (!instruction_D[20] & (Mux411))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux41~19_combout ),
	.datad(\REGISTER_FILE|Mux41~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~18 .lut_mask = 16'hFA50;
defparam \rdata2_EX~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N14
cycloneive_lcell_comb \rdata2_EX~19 (
// Equation(s):
// \rdata2_EX~19_combout  = (\always2~2_combout  & ((\rdata2_EX~18_combout ))) # (!\always2~2_combout  & (\portB~44_combout ))

	.dataa(\portB~44_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~18_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~19_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~19 .lut_mask = 16'hFA0A;
defparam \rdata2_EX~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N15
dffeas \rdata2_EX[22] (
	.clk(CLK),
	.d(\rdata2_EX~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[22]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[22] .is_wysiwyg = "true";
defparam \rdata2_EX[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N8
cycloneive_lcell_comb \rdata2_M~46 (
// Equation(s):
// \rdata2_M~46_combout  = (\rdata2_M[16]~1_combout  & ((\sw_forwarding_output~9_combout ) # ((\rdata2_M[16]~0_combout )))) # (!\rdata2_M[16]~1_combout  & (((rdata2_EX[22] & !\rdata2_M[16]~0_combout ))))

	.dataa(\sw_forwarding_output~9_combout ),
	.datab(rdata2_EX[22]),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\rdata2_M[16]~0_combout ),
	.cin(gnd),
	.combout(\rdata2_M~46_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~46 .lut_mask = 16'hF0AC;
defparam \rdata2_M~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N24
cycloneive_lcell_comb \imm_M~9 (
// Equation(s):
// \imm_M~9_combout  = (imm_EX[6] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(imm_EX[6]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\imm_M~9_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~9 .lut_mask = 16'h00CC;
defparam \imm_M~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N25
dffeas \imm_M[6] (
	.clk(CLK),
	.d(\imm_M~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[6]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[6] .is_wysiwyg = "true";
defparam \imm_M[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N28
cycloneive_lcell_comb \imm_WB[6]~feeder (
// Equation(s):
// \imm_WB[6]~feeder_combout  = imm_M[6]

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(imm_M[6]),
	.cin(gnd),
	.combout(\imm_WB[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \imm_WB[6]~feeder .lut_mask = 16'hFF00;
defparam \imm_WB[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N29
dffeas \imm_WB[6] (
	.clk(CLK),
	.d(\imm_WB[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[6]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[6] .is_wysiwyg = "true";
defparam \imm_WB[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N31
dffeas \dmemload_WB[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_22),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[22]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[22] .is_wysiwyg = "true";
defparam \dmemload_WB[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N6
cycloneive_lcell_comb \pc_plus_4_M~23 (
// Equation(s):
// \pc_plus_4_M~23_combout  = (pc_plus_4_EX[22] & !\wsel_M~0_combout )

	.dataa(pc_plus_4_EX[22]),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pc_plus_4_M~23_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~23 .lut_mask = 16'h0A0A;
defparam \pc_plus_4_M~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N7
dffeas \pc_plus_4_M[22] (
	.clk(CLK),
	.d(\pc_plus_4_M~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[22]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[22] .is_wysiwyg = "true";
defparam \pc_plus_4_M[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N10
cycloneive_lcell_comb \pc_plus_4_WB[22]~feeder (
// Equation(s):
// \pc_plus_4_WB[22]~feeder_combout  = pc_plus_4_M[22]

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pc_plus_4_M[22]),
	.cin(gnd),
	.combout(\pc_plus_4_WB[22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_WB[22]~feeder .lut_mask = 16'hFF00;
defparam \pc_plus_4_WB[22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N11
dffeas \pc_plus_4_WB[22] (
	.clk(CLK),
	.d(\pc_plus_4_WB[22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[22]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[22] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N21
dffeas \porto_WB[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_22),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[22]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[22] .is_wysiwyg = "true";
defparam \porto_WB[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N20
cycloneive_lcell_comb \wdat_WB[22]~20 (
// Equation(s):
// \wdat_WB[22]~20_combout  = (\wdat_WB[28]~0_combout  & ((pc_plus_4_WB[22]) # ((\wdat_WB[28]~1_combout )))) # (!\wdat_WB[28]~0_combout  & (((porto_WB[22] & !\wdat_WB[28]~1_combout ))))

	.dataa(\wdat_WB[28]~0_combout ),
	.datab(pc_plus_4_WB[22]),
	.datac(porto_WB[22]),
	.datad(\wdat_WB[28]~1_combout ),
	.cin(gnd),
	.combout(\wdat_WB[22]~20_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[22]~20 .lut_mask = 16'hAAD8;
defparam \wdat_WB[22]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N30
cycloneive_lcell_comb \wdat_WB[22]~21 (
// Equation(s):
// \wdat_WB[22]~21_combout  = (\wdat_WB[28]~1_combout  & ((\wdat_WB[22]~20_combout  & (imm_WB[6])) # (!\wdat_WB[22]~20_combout  & ((dmemload_WB[22]))))) # (!\wdat_WB[28]~1_combout  & (((\wdat_WB[22]~20_combout ))))

	.dataa(\wdat_WB[28]~1_combout ),
	.datab(imm_WB[6]),
	.datac(dmemload_WB[22]),
	.datad(\wdat_WB[22]~20_combout ),
	.cin(gnd),
	.combout(\wdat_WB[22]~21_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[22]~21 .lut_mask = 16'hDDA0;
defparam \wdat_WB[22]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N10
cycloneive_lcell_comb \rdata2_M~47 (
// Equation(s):
// \rdata2_M~47_combout  = (\rdata2_M~46_combout  & (((\wdat_WB[22]~21_combout )) # (!\rdata2_M[16]~0_combout ))) # (!\rdata2_M~46_combout  & (\rdata2_M[16]~0_combout  & ((ramiframload_22))))

	.dataa(\rdata2_M~46_combout ),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\wdat_WB[22]~21_combout ),
	.datad(ramiframload_22),
	.cin(gnd),
	.combout(\rdata2_M~47_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~47 .lut_mask = 16'hE6A2;
defparam \rdata2_M~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N4
cycloneive_lcell_comb \instruction_D~94 (
// Equation(s):
// \instruction_D~94_combout  = (\branch_or_jump~1_combout  & (iwait & ramiframload_7))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(iwait),
	.datad(ramiframload_7),
	.cin(gnd),
	.combout(\instruction_D~94_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~94 .lut_mask = 16'hA000;
defparam \instruction_D~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N5
dffeas \instruction_D[7] (
	.clk(CLK),
	.d(\instruction_D~94_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[7]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[7] .is_wysiwyg = "true";
defparam \instruction_D[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N10
cycloneive_lcell_comb \imm_EX~8 (
// Equation(s):
// \imm_EX~8_combout  = (\branch_or_jump~2_combout  & (instruction_D[7] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(instruction_D[7]),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\imm_EX~8_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~8 .lut_mask = 16'h8008;
defparam \imm_EX~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N5
dffeas \imm_EX[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\imm_EX~8_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[7]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[7] .is_wysiwyg = "true";
defparam \imm_EX[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N20
cycloneive_lcell_comb \imm_M~8 (
// Equation(s):
// \imm_M~8_combout  = (!\wsel_M~0_combout  & imm_EX[7])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(imm_EX[7]),
	.cin(gnd),
	.combout(\imm_M~8_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~8 .lut_mask = 16'h0F00;
defparam \imm_M~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y32_N21
dffeas \imm_M[7] (
	.clk(CLK),
	.d(\imm_M~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[7]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[7] .is_wysiwyg = "true";
defparam \imm_M[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N10
cycloneive_lcell_comb \sw_forwarding_output~8 (
// Equation(s):
// \sw_forwarding_output~8_combout  = (\lui_M~q  & (imm_M[7])) # (!\lui_M~q  & ((porto_M_23)))

	.dataa(\lui_M~q ),
	.datab(gnd),
	.datac(imm_M[7]),
	.datad(porto_M_23),
	.cin(gnd),
	.combout(\sw_forwarding_output~8_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~8 .lut_mask = 16'hF5A0;
defparam \sw_forwarding_output~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y29_N11
dffeas \imm_WB[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[7]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[7]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[7] .is_wysiwyg = "true";
defparam \imm_WB[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N12
cycloneive_lcell_comb \pc_plus_4[23]~42 (
// Equation(s):
// \pc_plus_4[23]~42_combout  = (pc_out_23 & (!\pc_plus_4[22]~41 )) # (!pc_out_23 & ((\pc_plus_4[22]~41 ) # (GND)))
// \pc_plus_4[23]~43  = CARRY((!\pc_plus_4[22]~41 ) # (!pc_out_23))

	.dataa(gnd),
	.datab(pc_out_23),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[22]~41 ),
	.combout(\pc_plus_4[23]~42_combout ),
	.cout(\pc_plus_4[23]~43 ));
// synopsys translate_off
defparam \pc_plus_4[23]~42 .lut_mask = 16'h3C3F;
defparam \pc_plus_4[23]~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N20
cycloneive_lcell_comb \pc_plus_4_D~22 (
// Equation(s):
// \pc_plus_4_D~22_combout  = (\pc_plus_4[23]~42_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(gnd),
	.datab(\branch_or_jump~1_combout ),
	.datac(iwait),
	.datad(\pc_plus_4[23]~42_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~22_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~22 .lut_mask = 16'hF300;
defparam \pc_plus_4_D~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N21
dffeas \pc_plus_4_D[23] (
	.clk(CLK),
	.d(\pc_plus_4_D~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[23]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[23] .is_wysiwyg = "true";
defparam \pc_plus_4_D[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N22
cycloneive_lcell_comb \pc_plus_4_EX~22 (
// Equation(s):
// \pc_plus_4_EX~22_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[23] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_D[23]),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~22_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~22 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N23
dffeas \pc_plus_4_EX[23] (
	.clk(CLK),
	.d(\pc_plus_4_EX~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[23]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[23] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N30
cycloneive_lcell_comb \pc_plus_4_M~22 (
// Equation(s):
// \pc_plus_4_M~22_combout  = (pc_plus_4_EX[23] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[23]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~22_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~22 .lut_mask = 16'h00CC;
defparam \pc_plus_4_M~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N31
dffeas \pc_plus_4_M[23] (
	.clk(CLK),
	.d(\pc_plus_4_M~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[23]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[23] .is_wysiwyg = "true";
defparam \pc_plus_4_M[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N17
dffeas \pc_plus_4_WB[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[23]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[23]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[23] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N25
dffeas \dmemload_WB[23] (
	.clk(CLK),
	.d(\dpif.dmemload [23]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[23]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[23] .is_wysiwyg = "true";
defparam \dmemload_WB[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N7
dffeas \porto_WB[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_23),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[23]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[23] .is_wysiwyg = "true";
defparam \porto_WB[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N6
cycloneive_lcell_comb \wdat_WB[23]~18 (
// Equation(s):
// \wdat_WB[23]~18_combout  = (\wdat_WB[28]~0_combout  & (((\wdat_WB[28]~1_combout )))) # (!\wdat_WB[28]~0_combout  & ((\wdat_WB[28]~1_combout  & (dmemload_WB[23])) # (!\wdat_WB[28]~1_combout  & ((porto_WB[23])))))

	.dataa(\wdat_WB[28]~0_combout ),
	.datab(dmemload_WB[23]),
	.datac(porto_WB[23]),
	.datad(\wdat_WB[28]~1_combout ),
	.cin(gnd),
	.combout(\wdat_WB[23]~18_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[23]~18 .lut_mask = 16'hEE50;
defparam \wdat_WB[23]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N16
cycloneive_lcell_comb \wdat_WB[23]~19 (
// Equation(s):
// \wdat_WB[23]~19_combout  = (\wdat_WB[28]~0_combout  & ((\wdat_WB[23]~18_combout  & (imm_WB[7])) # (!\wdat_WB[23]~18_combout  & ((pc_plus_4_WB[23]))))) # (!\wdat_WB[28]~0_combout  & (((\wdat_WB[23]~18_combout ))))

	.dataa(\wdat_WB[28]~0_combout ),
	.datab(imm_WB[7]),
	.datac(pc_plus_4_WB[23]),
	.datad(\wdat_WB[23]~18_combout ),
	.cin(gnd),
	.combout(\wdat_WB[23]~19_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[23]~19 .lut_mask = 16'hDDA0;
defparam \wdat_WB[23]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N20
cycloneive_lcell_comb \rdata2_EX~16 (
// Equation(s):
// \rdata2_EX~16_combout  = (instruction_D[20] & (Mux40)) # (!instruction_D[20] & ((Mux401)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux40~9_combout ),
	.datad(\REGISTER_FILE|Mux40~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~16 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N22
cycloneive_lcell_comb \rdata2_EX~17 (
// Equation(s):
// \rdata2_EX~17_combout  = (\always2~2_combout  & ((\rdata2_EX~16_combout ))) # (!\always2~2_combout  & (\portB~41_combout ))

	.dataa(\portB~41_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~16_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~17_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~17 .lut_mask = 16'hFA0A;
defparam \rdata2_EX~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N23
dffeas \rdata2_EX[23] (
	.clk(CLK),
	.d(\rdata2_EX~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[23]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[23] .is_wysiwyg = "true";
defparam \rdata2_EX[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N12
cycloneive_lcell_comb \rdata2_M~48 (
// Equation(s):
// \rdata2_M~48_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout ) # (ramiframload_23)))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[23] & (!\rdata2_M[16]~1_combout )))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(rdata2_EX[23]),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\dpif.dmemload [23]),
	.cin(gnd),
	.combout(\rdata2_M~48_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~48 .lut_mask = 16'hAEA4;
defparam \rdata2_M~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N24
cycloneive_lcell_comb \rdata2_M~49 (
// Equation(s):
// \rdata2_M~49_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~48_combout  & ((\wdat_WB[23]~19_combout ))) # (!\rdata2_M~48_combout  & (\sw_forwarding_output~8_combout )))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~48_combout ))))

	.dataa(\sw_forwarding_output~8_combout ),
	.datab(\wdat_WB[23]~19_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\rdata2_M~48_combout ),
	.cin(gnd),
	.combout(\rdata2_M~49_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~49 .lut_mask = 16'hCFA0;
defparam \rdata2_M~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N12
cycloneive_lcell_comb \imm_M~7 (
// Equation(s):
// \imm_M~7_combout  = (imm_EX[8] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(imm_EX[8]),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\imm_M~7_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~7 .lut_mask = 16'h0C0C;
defparam \imm_M~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N13
dffeas \imm_M[8] (
	.clk(CLK),
	.d(\imm_M~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[8]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[8] .is_wysiwyg = "true";
defparam \imm_M[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N25
dffeas \imm_WB[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[8]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[8]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[8] .is_wysiwyg = "true";
defparam \imm_WB[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N31
dffeas \dmemload_WB[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramiframload_24),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[24]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[24] .is_wysiwyg = "true";
defparam \dmemload_WB[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N26
cycloneive_lcell_comb \pc_plus_4_EX~25 (
// Equation(s):
// \pc_plus_4_EX~25_combout  = (pc_plus_4_D[24] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[24]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~25_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~25 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N27
dffeas \pc_plus_4_EX[24] (
	.clk(CLK),
	.d(\pc_plus_4_EX~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[24]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[24] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N14
cycloneive_lcell_comb \pc_plus_4_M~25 (
// Equation(s):
// \pc_plus_4_M~25_combout  = (pc_plus_4_EX[24] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(pc_plus_4_EX[24]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~25_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~25 .lut_mask = 16'h00CC;
defparam \pc_plus_4_M~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N15
dffeas \pc_plus_4_M[24] (
	.clk(CLK),
	.d(\pc_plus_4_M~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[24]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[24] .is_wysiwyg = "true";
defparam \pc_plus_4_M[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N13
dffeas \pc_plus_4_WB[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[24]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[24]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[24] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N3
dffeas \porto_WB[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_24),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[24]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[24] .is_wysiwyg = "true";
defparam \porto_WB[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N2
cycloneive_lcell_comb \wdat_WB[24]~16 (
// Equation(s):
// \wdat_WB[24]~16_combout  = (\wdat_WB[28]~0_combout  & ((pc_plus_4_WB[24]) # ((\wdat_WB[28]~1_combout )))) # (!\wdat_WB[28]~0_combout  & (((porto_WB[24] & !\wdat_WB[28]~1_combout ))))

	.dataa(\wdat_WB[28]~0_combout ),
	.datab(pc_plus_4_WB[24]),
	.datac(porto_WB[24]),
	.datad(\wdat_WB[28]~1_combout ),
	.cin(gnd),
	.combout(\wdat_WB[24]~16_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[24]~16 .lut_mask = 16'hAAD8;
defparam \wdat_WB[24]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N30
cycloneive_lcell_comb \wdat_WB[24]~17 (
// Equation(s):
// \wdat_WB[24]~17_combout  = (\wdat_WB[28]~1_combout  & ((\wdat_WB[24]~16_combout  & (imm_WB[8])) # (!\wdat_WB[24]~16_combout  & ((dmemload_WB[24]))))) # (!\wdat_WB[28]~1_combout  & (((\wdat_WB[24]~16_combout ))))

	.dataa(\wdat_WB[28]~1_combout ),
	.datab(imm_WB[8]),
	.datac(dmemload_WB[24]),
	.datad(\wdat_WB[24]~16_combout ),
	.cin(gnd),
	.combout(\wdat_WB[24]~17_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[24]~17 .lut_mask = 16'hDDA0;
defparam \wdat_WB[24]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N26
cycloneive_lcell_comb \rdata2_EX~14 (
// Equation(s):
// \rdata2_EX~14_combout  = (instruction_D[20] & (Mux39)) # (!instruction_D[20] & ((Mux391)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux39~9_combout ),
	.datad(\REGISTER_FILE|Mux39~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~14 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N8
cycloneive_lcell_comb \rdata2_EX~15 (
// Equation(s):
// \rdata2_EX~15_combout  = (\always2~2_combout  & ((\rdata2_EX~14_combout ))) # (!\always2~2_combout  & (\portB~38_combout ))

	.dataa(\portB~38_combout ),
	.datab(\always2~2_combout ),
	.datac(\rdata2_EX~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdata2_EX~15_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~15 .lut_mask = 16'hE2E2;
defparam \rdata2_EX~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N9
dffeas \rdata2_EX[24] (
	.clk(CLK),
	.d(\rdata2_EX~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[24]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[24] .is_wysiwyg = "true";
defparam \rdata2_EX[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N18
cycloneive_lcell_comb \sw_forwarding_output~7 (
// Equation(s):
// \sw_forwarding_output~7_combout  = (\lui_M~q  & (imm_M[8])) # (!\lui_M~q  & ((porto_M_24)))

	.dataa(gnd),
	.datab(\lui_M~q ),
	.datac(imm_M[8]),
	.datad(porto_M_24),
	.cin(gnd),
	.combout(\sw_forwarding_output~7_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~7 .lut_mask = 16'hF3C0;
defparam \sw_forwarding_output~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N28
cycloneive_lcell_comb \rdata2_M~50 (
// Equation(s):
// \rdata2_M~50_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & ((\rdata2_M[16]~1_combout  & ((\sw_forwarding_output~7_combout ))) # (!\rdata2_M[16]~1_combout  & (rdata2_EX[24]))))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(rdata2_EX[24]),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\sw_forwarding_output~7_combout ),
	.cin(gnd),
	.combout(\rdata2_M~50_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~50 .lut_mask = 16'hF4A4;
defparam \rdata2_M~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N14
cycloneive_lcell_comb \rdata2_M~51 (
// Equation(s):
// \rdata2_M~51_combout  = (\rdata2_M~50_combout  & ((\wdat_WB[24]~17_combout ) # ((!\rdata2_M[16]~0_combout )))) # (!\rdata2_M~50_combout  & (((\rdata2_M[16]~0_combout  & ramiframload_24))))

	.dataa(\wdat_WB[24]~17_combout ),
	.datab(\rdata2_M~50_combout ),
	.datac(\rdata2_M[16]~0_combout ),
	.datad(ramiframload_24),
	.cin(gnd),
	.combout(\rdata2_M~51_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~51 .lut_mask = 16'hBC8C;
defparam \rdata2_M~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N12
cycloneive_lcell_comb \imm_M~6 (
// Equation(s):
// \imm_M~6_combout  = (!\wsel_M~0_combout  & imm_EX[9])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(imm_EX[9]),
	.cin(gnd),
	.combout(\imm_M~6_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~6 .lut_mask = 16'h0F00;
defparam \imm_M~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N3
dffeas \imm_M[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\imm_M~6_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[9]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[9] .is_wysiwyg = "true";
defparam \imm_M[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N28
cycloneive_lcell_comb \imm_WB[9]~feeder (
// Equation(s):
// \imm_WB[9]~feeder_combout  = imm_M[9]

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(imm_M[9]),
	.cin(gnd),
	.combout(\imm_WB[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \imm_WB[9]~feeder .lut_mask = 16'hFF00;
defparam \imm_WB[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N29
dffeas \imm_WB[9] (
	.clk(CLK),
	.d(\imm_WB[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[9]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[9] .is_wysiwyg = "true";
defparam \imm_WB[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N16
cycloneive_lcell_comb \pc_plus_4[25]~46 (
// Equation(s):
// \pc_plus_4[25]~46_combout  = (pc_out_25 & (!\pc_plus_4[24]~45 )) # (!pc_out_25 & ((\pc_plus_4[24]~45 ) # (GND)))
// \pc_plus_4[25]~47  = CARRY((!\pc_plus_4[24]~45 ) # (!pc_out_25))

	.dataa(gnd),
	.datab(pc_out_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[24]~45 ),
	.combout(\pc_plus_4[25]~46_combout ),
	.cout(\pc_plus_4[25]~47 ));
// synopsys translate_off
defparam \pc_plus_4[25]~46 .lut_mask = 16'h3C3F;
defparam \pc_plus_4[25]~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N0
cycloneive_lcell_comb \pc_plus_4_D~24 (
// Equation(s):
// \pc_plus_4_D~24_combout  = (\pc_plus_4[25]~46_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(\pc_plus_4[25]~46_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\pc_plus_4_D~24_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~24 .lut_mask = 16'hF050;
defparam \pc_plus_4_D~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N1
dffeas \pc_plus_4_D[25] (
	.clk(CLK),
	.d(\pc_plus_4_D~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[25]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[25] .is_wysiwyg = "true";
defparam \pc_plus_4_D[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N16
cycloneive_lcell_comb \pc_plus_4_EX~24 (
// Equation(s):
// \pc_plus_4_EX~24_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[25] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_D[25]),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~24_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~24 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N17
dffeas \pc_plus_4_EX[25] (
	.clk(CLK),
	.d(\pc_plus_4_EX~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[25]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[25] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N30
cycloneive_lcell_comb \pc_plus_4_M~24 (
// Equation(s):
// \pc_plus_4_M~24_combout  = (pc_plus_4_EX[25] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_plus_4_EX[25]),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~24_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~24 .lut_mask = 16'h00F0;
defparam \pc_plus_4_M~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y39_N31
dffeas \pc_plus_4_M[25] (
	.clk(CLK),
	.d(\pc_plus_4_M~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[25]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[25] .is_wysiwyg = "true";
defparam \pc_plus_4_M[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N25
dffeas \pc_plus_4_WB[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[25]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[25]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[25] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N9
dffeas \dmemload_WB[25] (
	.clk(CLK),
	.d(\dpif.dmemload [25]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[25]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[25] .is_wysiwyg = "true";
defparam \dmemload_WB[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N3
dffeas \porto_WB[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_25),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[25]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[25] .is_wysiwyg = "true";
defparam \porto_WB[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N2
cycloneive_lcell_comb \wdat_WB[25]~14 (
// Equation(s):
// \wdat_WB[25]~14_combout  = (\wdat_WB[28]~0_combout  & (((\wdat_WB[28]~1_combout )))) # (!\wdat_WB[28]~0_combout  & ((\wdat_WB[28]~1_combout  & (dmemload_WB[25])) # (!\wdat_WB[28]~1_combout  & ((porto_WB[25])))))

	.dataa(\wdat_WB[28]~0_combout ),
	.datab(dmemload_WB[25]),
	.datac(porto_WB[25]),
	.datad(\wdat_WB[28]~1_combout ),
	.cin(gnd),
	.combout(\wdat_WB[25]~14_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[25]~14 .lut_mask = 16'hEE50;
defparam \wdat_WB[25]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N24
cycloneive_lcell_comb \wdat_WB[25]~15 (
// Equation(s):
// \wdat_WB[25]~15_combout  = (\wdat_WB[28]~0_combout  & ((\wdat_WB[25]~14_combout  & (imm_WB[9])) # (!\wdat_WB[25]~14_combout  & ((pc_plus_4_WB[25]))))) # (!\wdat_WB[28]~0_combout  & (((\wdat_WB[25]~14_combout ))))

	.dataa(\wdat_WB[28]~0_combout ),
	.datab(imm_WB[9]),
	.datac(pc_plus_4_WB[25]),
	.datad(\wdat_WB[25]~14_combout ),
	.cin(gnd),
	.combout(\wdat_WB[25]~15_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[25]~15 .lut_mask = 16'hDDA0;
defparam \wdat_WB[25]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N26
cycloneive_lcell_comb \sw_forwarding_output~6 (
// Equation(s):
// \sw_forwarding_output~6_combout  = (\lui_M~q  & (imm_M[9])) # (!\lui_M~q  & ((porto_M_25)))

	.dataa(imm_M[9]),
	.datab(gnd),
	.datac(porto_M_25),
	.datad(\lui_M~q ),
	.cin(gnd),
	.combout(\sw_forwarding_output~6_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~6 .lut_mask = 16'hAAF0;
defparam \sw_forwarding_output~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N30
cycloneive_lcell_comb \rdata2_M~52 (
// Equation(s):
// \rdata2_M~52_combout  = (\rdata2_M[16]~1_combout  & (((\rdata2_M[16]~0_combout )))) # (!\rdata2_M[16]~1_combout  & ((\rdata2_M[16]~0_combout  & ((ramiframload_25))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[25]))))

	.dataa(rdata2_EX[25]),
	.datab(\rdata2_M[16]~1_combout ),
	.datac(\dpif.dmemload [25]),
	.datad(\rdata2_M[16]~0_combout ),
	.cin(gnd),
	.combout(\rdata2_M~52_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~52 .lut_mask = 16'hFC22;
defparam \rdata2_M~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N12
cycloneive_lcell_comb \rdata2_M~53 (
// Equation(s):
// \rdata2_M~53_combout  = (\rdata2_M~52_combout  & ((\wdat_WB[25]~15_combout ) # ((!\rdata2_M[16]~1_combout )))) # (!\rdata2_M~52_combout  & (((\sw_forwarding_output~6_combout  & \rdata2_M[16]~1_combout ))))

	.dataa(\wdat_WB[25]~15_combout ),
	.datab(\sw_forwarding_output~6_combout ),
	.datac(\rdata2_M~52_combout ),
	.datad(\rdata2_M[16]~1_combout ),
	.cin(gnd),
	.combout(\rdata2_M~53_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~53 .lut_mask = 16'hACF0;
defparam \rdata2_M~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N29
dffeas \dmemload_WB[26] (
	.clk(CLK),
	.d(\dpif.dmemload [26]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[26]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[26] .is_wysiwyg = "true";
defparam \dmemload_WB[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N0
cycloneive_lcell_comb \imm_M~5 (
// Equation(s):
// \imm_M~5_combout  = (!\wsel_M~0_combout  & imm_EX[10])

	.dataa(\wsel_M~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(imm_EX[10]),
	.cin(gnd),
	.combout(\imm_M~5_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~5 .lut_mask = 16'h5500;
defparam \imm_M~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N1
dffeas \imm_M[10] (
	.clk(CLK),
	.d(\imm_M~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[10]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[10] .is_wysiwyg = "true";
defparam \imm_M[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N5
dffeas \imm_WB[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[10]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[10]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[10] .is_wysiwyg = "true";
defparam \imm_WB[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N28
cycloneive_lcell_comb \pc_plus_4_EX~27 (
// Equation(s):
// \pc_plus_4_EX~27_combout  = (pc_plus_4_D[26] & (\branch_or_jump~2_combout  & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(pc_plus_4_D[26]),
	.datab(\branch_taken~0_combout ),
	.datac(\branch_or_jump~2_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~27_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~27 .lut_mask = 16'h8020;
defparam \pc_plus_4_EX~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N29
dffeas \pc_plus_4_EX[26] (
	.clk(CLK),
	.d(\pc_plus_4_EX~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[26]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[26] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N14
cycloneive_lcell_comb \pc_plus_4_M~27 (
// Equation(s):
// \pc_plus_4_M~27_combout  = (!\wsel_M~0_combout  & pc_plus_4_EX[26])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(pc_plus_4_EX[26]),
	.cin(gnd),
	.combout(\pc_plus_4_M~27_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~27 .lut_mask = 16'h0F00;
defparam \pc_plus_4_M~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N15
dffeas \pc_plus_4_M[26] (
	.clk(CLK),
	.d(\pc_plus_4_M~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[26]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[26] .is_wysiwyg = "true";
defparam \pc_plus_4_M[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N17
dffeas \pc_plus_4_WB[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[26]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[26]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[26] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N3
dffeas \porto_WB[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_26),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[26]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[26] .is_wysiwyg = "true";
defparam \porto_WB[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N2
cycloneive_lcell_comb \wdat_WB[26]~12 (
// Equation(s):
// \wdat_WB[26]~12_combout  = (\wdat_WB[28]~0_combout  & ((pc_plus_4_WB[26]) # ((\wdat_WB[28]~1_combout )))) # (!\wdat_WB[28]~0_combout  & (((porto_WB[26] & !\wdat_WB[28]~1_combout ))))

	.dataa(\wdat_WB[28]~0_combout ),
	.datab(pc_plus_4_WB[26]),
	.datac(porto_WB[26]),
	.datad(\wdat_WB[28]~1_combout ),
	.cin(gnd),
	.combout(\wdat_WB[26]~12_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[26]~12 .lut_mask = 16'hAAD8;
defparam \wdat_WB[26]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N4
cycloneive_lcell_comb \wdat_WB[26]~13 (
// Equation(s):
// \wdat_WB[26]~13_combout  = (\wdat_WB[28]~1_combout  & ((\wdat_WB[26]~12_combout  & ((imm_WB[10]))) # (!\wdat_WB[26]~12_combout  & (dmemload_WB[26])))) # (!\wdat_WB[28]~1_combout  & (((\wdat_WB[26]~12_combout ))))

	.dataa(\wdat_WB[28]~1_combout ),
	.datab(dmemload_WB[26]),
	.datac(imm_WB[10]),
	.datad(\wdat_WB[26]~12_combout ),
	.cin(gnd),
	.combout(\wdat_WB[26]~13_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[26]~13 .lut_mask = 16'hF588;
defparam \wdat_WB[26]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N10
cycloneive_lcell_comb \portB~30 (
// Equation(s):
// \portB~30_combout  = (\Equal3~2_combout  & (((\portB~14_combout )))) # (!\Equal3~2_combout  & ((\portB~14_combout  & ((\sign_ext[16]~0_combout ))) # (!\portB~14_combout  & (rdata2_EX[26]))))

	.dataa(rdata2_EX[26]),
	.datab(\sign_ext[16]~0_combout ),
	.datac(\Equal3~2_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~30_combout ),
	.cout());
// synopsys translate_off
defparam \portB~30 .lut_mask = 16'hFC0A;
defparam \portB~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N6
cycloneive_lcell_comb \portB~31 (
// Equation(s):
// \portB~31_combout  = (\Equal3~2_combout  & ((\portB~30_combout  & (\sw_forwarding_output~5_combout )) # (!\portB~30_combout  & ((\wdat_WB[26]~13_combout ))))) # (!\Equal3~2_combout  & (((\portB~30_combout ))))

	.dataa(\sw_forwarding_output~5_combout ),
	.datab(\wdat_WB[26]~13_combout ),
	.datac(\Equal3~2_combout ),
	.datad(\portB~30_combout ),
	.cin(gnd),
	.combout(\portB~31_combout ),
	.cout());
// synopsys translate_off
defparam \portB~31 .lut_mask = 16'hAFC0;
defparam \portB~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N20
cycloneive_lcell_comb \portB~32 (
// Equation(s):
// \portB~32_combout  = (\portB~31_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(gnd),
	.datab(\ShiftOp_EX~q ),
	.datac(\Equal3~2_combout ),
	.datad(\portB~31_combout ),
	.cin(gnd),
	.combout(\portB~32_combout ),
	.cout());
// synopsys translate_off
defparam \portB~32 .lut_mask = 16'hF300;
defparam \portB~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N2
cycloneive_lcell_comb \rdata2_EX~10 (
// Equation(s):
// \rdata2_EX~10_combout  = (instruction_D[20] & ((Mux37))) # (!instruction_D[20] & (Mux371))

	.dataa(gnd),
	.datab(instruction_D[20]),
	.datac(\REGISTER_FILE|Mux37~19_combout ),
	.datad(\REGISTER_FILE|Mux37~9_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~10 .lut_mask = 16'hFC30;
defparam \rdata2_EX~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N20
cycloneive_lcell_comb \rdata2_EX~11 (
// Equation(s):
// \rdata2_EX~11_combout  = (\always2~2_combout  & ((\rdata2_EX~10_combout ))) # (!\always2~2_combout  & (\portB~32_combout ))

	.dataa(gnd),
	.datab(\portB~32_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~10_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~11_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~11 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N21
dffeas \rdata2_EX[26] (
	.clk(CLK),
	.d(\rdata2_EX~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[26]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[26] .is_wysiwyg = "true";
defparam \rdata2_EX[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N14
cycloneive_lcell_comb \rdata2_M~54 (
// Equation(s):
// \rdata2_M~54_combout  = (\rdata2_M[16]~1_combout  & ((\sw_forwarding_output~5_combout ) # ((\rdata2_M[16]~0_combout )))) # (!\rdata2_M[16]~1_combout  & (((rdata2_EX[26] & !\rdata2_M[16]~0_combout ))))

	.dataa(\sw_forwarding_output~5_combout ),
	.datab(rdata2_EX[26]),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\rdata2_M[16]~0_combout ),
	.cin(gnd),
	.combout(\rdata2_M~54_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~54 .lut_mask = 16'hF0AC;
defparam \rdata2_M~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N6
cycloneive_lcell_comb \rdata2_M~55 (
// Equation(s):
// \rdata2_M~55_combout  = (\rdata2_M[16]~0_combout  & ((\rdata2_M~54_combout  & (\wdat_WB[26]~13_combout )) # (!\rdata2_M~54_combout  & ((ramiframload_26))))) # (!\rdata2_M[16]~0_combout  & (((\rdata2_M~54_combout ))))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(\wdat_WB[26]~13_combout ),
	.datac(\rdata2_M~54_combout ),
	.datad(\dpif.dmemload [26]),
	.cin(gnd),
	.combout(\rdata2_M~55_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~55 .lut_mask = 16'hDAD0;
defparam \rdata2_M~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N20
cycloneive_lcell_comb \pc_plus_4[27]~50 (
// Equation(s):
// \pc_plus_4[27]~50_combout  = (pc_out_27 & (!\pc_plus_4[26]~49 )) # (!pc_out_27 & ((\pc_plus_4[26]~49 ) # (GND)))
// \pc_plus_4[27]~51  = CARRY((!\pc_plus_4[26]~49 ) # (!pc_out_27))

	.dataa(pc_out_27),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\pc_plus_4[26]~49 ),
	.combout(\pc_plus_4[27]~50_combout ),
	.cout(\pc_plus_4[27]~51 ));
// synopsys translate_off
defparam \pc_plus_4[27]~50 .lut_mask = 16'h5A5F;
defparam \pc_plus_4[27]~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N8
cycloneive_lcell_comb \pc_plus_4_D~26 (
// Equation(s):
// \pc_plus_4_D~26_combout  = (\pc_plus_4[27]~50_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(\branch_or_jump~1_combout ),
	.datab(gnd),
	.datac(\pc_plus_4[27]~50_combout ),
	.datad(iwait),
	.cin(gnd),
	.combout(\pc_plus_4_D~26_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~26 .lut_mask = 16'hF050;
defparam \pc_plus_4_D~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N9
dffeas \pc_plus_4_D[27] (
	.clk(CLK),
	.d(\pc_plus_4_D~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[27]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[27] .is_wysiwyg = "true";
defparam \pc_plus_4_D[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N24
cycloneive_lcell_comb \pc_plus_4_EX~26 (
// Equation(s):
// \pc_plus_4_EX~26_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[27] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(\predicted_M~q ),
	.datac(pc_plus_4_D[27]),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~26_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~26 .lut_mask = 16'h8020;
defparam \pc_plus_4_EX~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N25
dffeas \pc_plus_4_EX[27] (
	.clk(CLK),
	.d(\pc_plus_4_EX~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[27]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[27] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N24
cycloneive_lcell_comb \pc_plus_4_M~26 (
// Equation(s):
// \pc_plus_4_M~26_combout  = (!\wsel_M~0_combout  & pc_plus_4_EX[27])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(pc_plus_4_EX[27]),
	.cin(gnd),
	.combout(\pc_plus_4_M~26_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~26 .lut_mask = 16'h0F00;
defparam \pc_plus_4_M~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N25
dffeas \pc_plus_4_M[27] (
	.clk(CLK),
	.d(\pc_plus_4_M~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[27]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[27] .is_wysiwyg = "true";
defparam \pc_plus_4_M[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N29
dffeas \pc_plus_4_WB[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[27]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[27]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[27] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N5
dffeas \porto_WB[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_27),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[27]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[27] .is_wysiwyg = "true";
defparam \porto_WB[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N4
cycloneive_lcell_comb \wdat_WB[27]~10 (
// Equation(s):
// \wdat_WB[27]~10_combout  = (\wdat_WB[28]~0_combout  & (((\wdat_WB[28]~1_combout )))) # (!\wdat_WB[28]~0_combout  & ((\wdat_WB[28]~1_combout  & (dmemload_WB[27])) # (!\wdat_WB[28]~1_combout  & ((porto_WB[27])))))

	.dataa(dmemload_WB[27]),
	.datab(\wdat_WB[28]~0_combout ),
	.datac(porto_WB[27]),
	.datad(\wdat_WB[28]~1_combout ),
	.cin(gnd),
	.combout(\wdat_WB[27]~10_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[27]~10 .lut_mask = 16'hEE30;
defparam \wdat_WB[27]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N28
cycloneive_lcell_comb \wdat_WB[27]~11 (
// Equation(s):
// \wdat_WB[27]~11_combout  = (\wdat_WB[28]~0_combout  & ((\wdat_WB[27]~10_combout  & (imm_WB[11])) # (!\wdat_WB[27]~10_combout  & ((pc_plus_4_WB[27]))))) # (!\wdat_WB[28]~0_combout  & (((\wdat_WB[27]~10_combout ))))

	.dataa(imm_WB[11]),
	.datab(\wdat_WB[28]~0_combout ),
	.datac(pc_plus_4_WB[27]),
	.datad(\wdat_WB[27]~10_combout ),
	.cin(gnd),
	.combout(\wdat_WB[27]~11_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[27]~11 .lut_mask = 16'hBBC0;
defparam \wdat_WB[27]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N30
cycloneive_lcell_comb \imm_M~4 (
// Equation(s):
// \imm_M~4_combout  = (imm_EX[11] & !\wsel_M~0_combout )

	.dataa(imm_EX[11]),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\imm_M~4_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~4 .lut_mask = 16'h0A0A;
defparam \imm_M~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N31
dffeas \imm_M[11] (
	.clk(CLK),
	.d(\imm_M~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[11]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[11] .is_wysiwyg = "true";
defparam \imm_M[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N2
cycloneive_lcell_comb \sw_forwarding_output~4 (
// Equation(s):
// \sw_forwarding_output~4_combout  = (\lui_M~q  & ((imm_M[11]))) # (!\lui_M~q  & (porto_M_27))

	.dataa(porto_M_27),
	.datab(\lui_M~q ),
	.datac(gnd),
	.datad(imm_M[11]),
	.cin(gnd),
	.combout(\sw_forwarding_output~4_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~4 .lut_mask = 16'hEE22;
defparam \sw_forwarding_output~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N14
cycloneive_lcell_comb \rdata2_M~56 (
// Equation(s):
// \rdata2_M~56_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout ) # (ramiframload_27)))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[27] & (!\rdata2_M[16]~1_combout )))

	.dataa(rdata2_EX[27]),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\dpif.dmemload [27]),
	.cin(gnd),
	.combout(\rdata2_M~56_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~56 .lut_mask = 16'hCEC2;
defparam \rdata2_M~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N0
cycloneive_lcell_comb \rdata2_M~57 (
// Equation(s):
// \rdata2_M~57_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~56_combout  & (\wdat_WB[27]~11_combout )) # (!\rdata2_M~56_combout  & ((\sw_forwarding_output~4_combout ))))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~56_combout ))))

	.dataa(\rdata2_M[16]~1_combout ),
	.datab(\wdat_WB[27]~11_combout ),
	.datac(\sw_forwarding_output~4_combout ),
	.datad(\rdata2_M~56_combout ),
	.cin(gnd),
	.combout(\rdata2_M~57_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~57 .lut_mask = 16'hDDA0;
defparam \rdata2_M~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N19
dffeas \porto_WB[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_28),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[28]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[28] .is_wysiwyg = "true";
defparam \porto_WB[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N18
cycloneive_lcell_comb \wdat_WB[28]~8 (
// Equation(s):
// \wdat_WB[28]~8_combout  = (\wdat_WB[28]~0_combout  & ((pc_plus_4_WB[28]) # ((\wdat_WB[28]~1_combout )))) # (!\wdat_WB[28]~0_combout  & (((porto_WB[28] & !\wdat_WB[28]~1_combout ))))

	.dataa(pc_plus_4_WB[28]),
	.datab(\wdat_WB[28]~0_combout ),
	.datac(porto_WB[28]),
	.datad(\wdat_WB[28]~1_combout ),
	.cin(gnd),
	.combout(\wdat_WB[28]~8_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[28]~8 .lut_mask = 16'hCCB8;
defparam \wdat_WB[28]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N2
cycloneive_lcell_comb \instruction_D~89 (
// Equation(s):
// \instruction_D~89_combout  = (iwait & (\branch_or_jump~1_combout  & ramiframload_12))

	.dataa(iwait),
	.datab(gnd),
	.datac(\branch_or_jump~1_combout ),
	.datad(\dpif.dmemload [12]),
	.cin(gnd),
	.combout(\instruction_D~89_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~89 .lut_mask = 16'hA000;
defparam \instruction_D~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N3
dffeas \instruction_D[12] (
	.clk(CLK),
	.d(\instruction_D~89_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[12]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[12] .is_wysiwyg = "true";
defparam \instruction_D[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N10
cycloneive_lcell_comb \imm_EX~3 (
// Equation(s):
// \imm_EX~3_combout  = (\branch_or_jump~2_combout  & (instruction_D[12] & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(instruction_D[12]),
	.datac(\branch_taken~0_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\imm_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~3 .lut_mask = 16'h8008;
defparam \imm_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N11
dffeas \imm_EX[12] (
	.clk(CLK),
	.d(\imm_EX~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[12]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[12] .is_wysiwyg = "true";
defparam \imm_EX[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N8
cycloneive_lcell_comb \imm_M~3 (
// Equation(s):
// \imm_M~3_combout  = (imm_EX[12] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(imm_EX[12]),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\imm_M~3_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~3 .lut_mask = 16'h00CC;
defparam \imm_M~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N9
dffeas \imm_M[12] (
	.clk(CLK),
	.d(\imm_M~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[12]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[12] .is_wysiwyg = "true";
defparam \imm_M[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N1
dffeas \imm_WB[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[12]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[12]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[12] .is_wysiwyg = "true";
defparam \imm_WB[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N0
cycloneive_lcell_comb \wdat_WB[28]~9 (
// Equation(s):
// \wdat_WB[28]~9_combout  = (\wdat_WB[28]~8_combout  & (((imm_WB[12]) # (!\wdat_WB[28]~1_combout )))) # (!\wdat_WB[28]~8_combout  & (dmemload_WB[28] & ((\wdat_WB[28]~1_combout ))))

	.dataa(dmemload_WB[28]),
	.datab(\wdat_WB[28]~8_combout ),
	.datac(imm_WB[12]),
	.datad(\wdat_WB[28]~1_combout ),
	.cin(gnd),
	.combout(\wdat_WB[28]~9_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[28]~9 .lut_mask = 16'hE2CC;
defparam \wdat_WB[28]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N26
cycloneive_lcell_comb \portB~24 (
// Equation(s):
// \portB~24_combout  = (\Equal3~2_combout  & (((\wdat_WB[28]~9_combout ) # (\portB~14_combout )))) # (!\Equal3~2_combout  & (rdata2_EX[28] & ((!\portB~14_combout ))))

	.dataa(rdata2_EX[28]),
	.datab(\wdat_WB[28]~9_combout ),
	.datac(\Equal3~2_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~24_combout ),
	.cout());
// synopsys translate_off
defparam \portB~24 .lut_mask = 16'hF0CA;
defparam \portB~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N10
cycloneive_lcell_comb \portB~25 (
// Equation(s):
// \portB~25_combout  = (\portB~14_combout  & ((\portB~24_combout  & (\sw_forwarding_output~3_combout )) # (!\portB~24_combout  & ((\sign_ext[16]~0_combout ))))) # (!\portB~14_combout  & (((\portB~24_combout ))))

	.dataa(\sw_forwarding_output~3_combout ),
	.datab(\sign_ext[16]~0_combout ),
	.datac(\portB~14_combout ),
	.datad(\portB~24_combout ),
	.cin(gnd),
	.combout(\portB~25_combout ),
	.cout());
// synopsys translate_off
defparam \portB~25 .lut_mask = 16'hAFC0;
defparam \portB~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N12
cycloneive_lcell_comb \portB~26 (
// Equation(s):
// \portB~26_combout  = (\portB~25_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(\ShiftOp_EX~q ),
	.datab(\Equal3~2_combout ),
	.datac(gnd),
	.datad(\portB~25_combout ),
	.cin(gnd),
	.combout(\portB~26_combout ),
	.cout());
// synopsys translate_off
defparam \portB~26 .lut_mask = 16'hDD00;
defparam \portB~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N6
cycloneive_lcell_comb \rdata2_EX~6 (
// Equation(s):
// \rdata2_EX~6_combout  = (instruction_D[20] & (Mux35)) # (!instruction_D[20] & ((Mux351)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux35~9_combout ),
	.datad(\REGISTER_FILE|Mux35~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~6 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N12
cycloneive_lcell_comb \rdata2_EX~7 (
// Equation(s):
// \rdata2_EX~7_combout  = (\always2~2_combout  & ((\rdata2_EX~6_combout ))) # (!\always2~2_combout  & (\portB~26_combout ))

	.dataa(gnd),
	.datab(\portB~26_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~6_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~7_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~7 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N13
dffeas \rdata2_EX[28] (
	.clk(CLK),
	.d(\rdata2_EX~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[28]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[28] .is_wysiwyg = "true";
defparam \rdata2_EX[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N18
cycloneive_lcell_comb \sw_forwarding_output~3 (
// Equation(s):
// \sw_forwarding_output~3_combout  = (\lui_M~q  & (imm_M[12])) # (!\lui_M~q  & ((porto_M_28)))

	.dataa(gnd),
	.datab(\lui_M~q ),
	.datac(imm_M[12]),
	.datad(porto_M_28),
	.cin(gnd),
	.combout(\sw_forwarding_output~3_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~3 .lut_mask = 16'hF3C0;
defparam \sw_forwarding_output~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N10
cycloneive_lcell_comb \rdata2_M~58 (
// Equation(s):
// \rdata2_M~58_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M[16]~0_combout ) # ((\sw_forwarding_output~3_combout )))) # (!\rdata2_M[16]~1_combout  & (!\rdata2_M[16]~0_combout  & (rdata2_EX[28])))

	.dataa(\rdata2_M[16]~1_combout ),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(rdata2_EX[28]),
	.datad(\sw_forwarding_output~3_combout ),
	.cin(gnd),
	.combout(\rdata2_M~58_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~58 .lut_mask = 16'hBA98;
defparam \rdata2_M~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N16
cycloneive_lcell_comb \rdata2_M~59 (
// Equation(s):
// \rdata2_M~59_combout  = (\rdata2_M[16]~0_combout  & ((\rdata2_M~58_combout  & (\wdat_WB[28]~9_combout )) # (!\rdata2_M~58_combout  & ((ramiframload_28))))) # (!\rdata2_M[16]~0_combout  & (((\rdata2_M~58_combout ))))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(\wdat_WB[28]~9_combout ),
	.datac(\dpif.dmemload [28]),
	.datad(\rdata2_M~58_combout ),
	.cin(gnd),
	.combout(\rdata2_M~59_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~59 .lut_mask = 16'hDDA0;
defparam \rdata2_M~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N2
cycloneive_lcell_comb \instruction_D~88 (
// Equation(s):
// \instruction_D~88_combout  = (iwait & (\branch_or_jump~1_combout  & ramiframload_13))

	.dataa(gnd),
	.datab(iwait),
	.datac(\branch_or_jump~1_combout ),
	.datad(\dpif.dmemload [13]),
	.cin(gnd),
	.combout(\instruction_D~88_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~88 .lut_mask = 16'hC000;
defparam \instruction_D~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N3
dffeas \instruction_D[13] (
	.clk(CLK),
	.d(\instruction_D~88_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[13]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[13] .is_wysiwyg = "true";
defparam \instruction_D[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N20
cycloneive_lcell_comb \imm_EX~2 (
// Equation(s):
// \imm_EX~2_combout  = (\branch_or_jump~2_combout  & (instruction_D[13] & (\branch_taken~0_combout  $ (!\predicted_M~q ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(instruction_D[13]),
	.datac(\branch_taken~0_combout ),
	.datad(\predicted_M~q ),
	.cin(gnd),
	.combout(\imm_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \imm_EX~2 .lut_mask = 16'h8008;
defparam \imm_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N21
dffeas \imm_EX[13] (
	.clk(CLK),
	.d(\imm_EX~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_EX[13]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_EX[13] .is_wysiwyg = "true";
defparam \imm_EX[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N16
cycloneive_lcell_comb \imm_M~2 (
// Equation(s):
// \imm_M~2_combout  = (!\wsel_M~0_combout  & imm_EX[13])

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(imm_EX[13]),
	.cin(gnd),
	.combout(\imm_M~2_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~2 .lut_mask = 16'h0F00;
defparam \imm_M~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y28_N17
dffeas \imm_M[13] (
	.clk(CLK),
	.d(\imm_M~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[13]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[13] .is_wysiwyg = "true";
defparam \imm_M[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N2
cycloneive_lcell_comb \sw_forwarding_output~2 (
// Equation(s):
// \sw_forwarding_output~2_combout  = (\lui_M~q  & (imm_M[13])) # (!\lui_M~q  & ((porto_M_29)))

	.dataa(gnd),
	.datab(imm_M[13]),
	.datac(\lui_M~q ),
	.datad(porto_M_29),
	.cin(gnd),
	.combout(\sw_forwarding_output~2_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~2 .lut_mask = 16'hCFC0;
defparam \sw_forwarding_output~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N4
cycloneive_lcell_comb \imm_WB[13]~feeder (
// Equation(s):
// \imm_WB[13]~feeder_combout  = imm_M[13]

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(imm_M[13]),
	.cin(gnd),
	.combout(\imm_WB[13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \imm_WB[13]~feeder .lut_mask = 16'hFF00;
defparam \imm_WB[13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N5
dffeas \imm_WB[13] (
	.clk(CLK),
	.d(\imm_WB[13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[13]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[13] .is_wysiwyg = "true";
defparam \imm_WB[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N10
cycloneive_lcell_comb \pc_plus_4_M~28 (
// Equation(s):
// \pc_plus_4_M~28_combout  = (pc_plus_4_EX[29] & !\wsel_M~0_combout )

	.dataa(pc_plus_4_EX[29]),
	.datab(gnd),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~28_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~28 .lut_mask = 16'h00AA;
defparam \pc_plus_4_M~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N11
dffeas \pc_plus_4_M[29] (
	.clk(CLK),
	.d(\pc_plus_4_M~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[29]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[29] .is_wysiwyg = "true";
defparam \pc_plus_4_M[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N13
dffeas \pc_plus_4_WB[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[29]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[29]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[29] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N1
dffeas \dmemload_WB[29] (
	.clk(CLK),
	.d(\dpif.dmemload [29]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[29]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[29] .is_wysiwyg = "true";
defparam \dmemload_WB[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N3
dffeas \porto_WB[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_29),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[29]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[29] .is_wysiwyg = "true";
defparam \porto_WB[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N2
cycloneive_lcell_comb \wdat_WB[29]~6 (
// Equation(s):
// \wdat_WB[29]~6_combout  = (\wdat_WB[28]~1_combout  & ((dmemload_WB[29]) # ((\wdat_WB[28]~0_combout )))) # (!\wdat_WB[28]~1_combout  & (((porto_WB[29] & !\wdat_WB[28]~0_combout ))))

	.dataa(\wdat_WB[28]~1_combout ),
	.datab(dmemload_WB[29]),
	.datac(porto_WB[29]),
	.datad(\wdat_WB[28]~0_combout ),
	.cin(gnd),
	.combout(\wdat_WB[29]~6_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[29]~6 .lut_mask = 16'hAAD8;
defparam \wdat_WB[29]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N12
cycloneive_lcell_comb \wdat_WB[29]~7 (
// Equation(s):
// \wdat_WB[29]~7_combout  = (\wdat_WB[28]~0_combout  & ((\wdat_WB[29]~6_combout  & (imm_WB[13])) # (!\wdat_WB[29]~6_combout  & ((pc_plus_4_WB[29]))))) # (!\wdat_WB[28]~0_combout  & (((\wdat_WB[29]~6_combout ))))

	.dataa(\wdat_WB[28]~0_combout ),
	.datab(imm_WB[13]),
	.datac(pc_plus_4_WB[29]),
	.datad(\wdat_WB[29]~6_combout ),
	.cin(gnd),
	.combout(\wdat_WB[29]~7_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[29]~7 .lut_mask = 16'hDDA0;
defparam \wdat_WB[29]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N18
cycloneive_lcell_comb \portB~21 (
// Equation(s):
// \portB~21_combout  = (\portB~14_combout  & (((\Equal3~2_combout )))) # (!\portB~14_combout  & ((\Equal3~2_combout  & (\wdat_WB[29]~7_combout )) # (!\Equal3~2_combout  & ((rdata2_EX[29])))))

	.dataa(\wdat_WB[29]~7_combout ),
	.datab(rdata2_EX[29]),
	.datac(\portB~14_combout ),
	.datad(\Equal3~2_combout ),
	.cin(gnd),
	.combout(\portB~21_combout ),
	.cout());
// synopsys translate_off
defparam \portB~21 .lut_mask = 16'hFA0C;
defparam \portB~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N28
cycloneive_lcell_comb \portB~22 (
// Equation(s):
// \portB~22_combout  = (\portB~14_combout  & ((\portB~21_combout  & ((\sw_forwarding_output~2_combout ))) # (!\portB~21_combout  & (\sign_ext[16]~0_combout )))) # (!\portB~14_combout  & (((\portB~21_combout ))))

	.dataa(\portB~14_combout ),
	.datab(\sign_ext[16]~0_combout ),
	.datac(\sw_forwarding_output~2_combout ),
	.datad(\portB~21_combout ),
	.cin(gnd),
	.combout(\portB~22_combout ),
	.cout());
// synopsys translate_off
defparam \portB~22 .lut_mask = 16'hF588;
defparam \portB~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N28
cycloneive_lcell_comb \portB~23 (
// Equation(s):
// \portB~23_combout  = (\portB~22_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(\ShiftOp_EX~q ),
	.datab(\Equal3~2_combout ),
	.datac(gnd),
	.datad(\portB~22_combout ),
	.cin(gnd),
	.combout(\portB~23_combout ),
	.cout());
// synopsys translate_off
defparam \portB~23 .lut_mask = 16'hDD00;
defparam \portB~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N0
cycloneive_lcell_comb \rdata2_EX~4 (
// Equation(s):
// \rdata2_EX~4_combout  = (instruction_D[20] & (Mux34)) # (!instruction_D[20] & ((Mux341)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux34~9_combout ),
	.datad(\REGISTER_FILE|Mux34~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~4 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N22
cycloneive_lcell_comb \rdata2_EX~5 (
// Equation(s):
// \rdata2_EX~5_combout  = (\always2~2_combout  & ((\rdata2_EX~4_combout ))) # (!\always2~2_combout  & (\portB~23_combout ))

	.dataa(gnd),
	.datab(\portB~23_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~4_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~5_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~5 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N23
dffeas \rdata2_EX[29] (
	.clk(CLK),
	.d(\rdata2_EX~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[29]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[29] .is_wysiwyg = "true";
defparam \rdata2_EX[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N6
cycloneive_lcell_comb \rdata2_M~60 (
// Equation(s):
// \rdata2_M~60_combout  = (\rdata2_M[16]~1_combout  & (\rdata2_M[16]~0_combout )) # (!\rdata2_M[16]~1_combout  & ((\rdata2_M[16]~0_combout  & ((ramiframload_29))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[29]))))

	.dataa(\rdata2_M[16]~1_combout ),
	.datab(\rdata2_M[16]~0_combout ),
	.datac(rdata2_EX[29]),
	.datad(\dpif.dmemload [29]),
	.cin(gnd),
	.combout(\rdata2_M~60_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~60 .lut_mask = 16'hDC98;
defparam \rdata2_M~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N0
cycloneive_lcell_comb \rdata2_M~61 (
// Equation(s):
// \rdata2_M~61_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~60_combout  & ((\wdat_WB[29]~7_combout ))) # (!\rdata2_M~60_combout  & (\sw_forwarding_output~2_combout )))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~60_combout ))))

	.dataa(\rdata2_M[16]~1_combout ),
	.datab(\sw_forwarding_output~2_combout ),
	.datac(\wdat_WB[29]~7_combout ),
	.datad(\rdata2_M~60_combout ),
	.cin(gnd),
	.combout(\rdata2_M~61_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~61 .lut_mask = 16'hF588;
defparam \rdata2_M~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N20
cycloneive_lcell_comb \imm_M~1 (
// Equation(s):
// \imm_M~1_combout  = (imm_EX[14] & !\wsel_M~0_combout )

	.dataa(imm_EX[14]),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\imm_M~1_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~1 .lut_mask = 16'h0A0A;
defparam \imm_M~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N21
dffeas \imm_M[14] (
	.clk(CLK),
	.d(\imm_M~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[14]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[14] .is_wysiwyg = "true";
defparam \imm_M[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N9
dffeas \imm_WB[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(imm_M[14]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[14]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[14] .is_wysiwyg = "true";
defparam \imm_WB[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y34_N21
dffeas \porto_WB[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_30),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[30]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[30] .is_wysiwyg = "true";
defparam \porto_WB[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N4
cycloneive_lcell_comb \pc_plus_4_D~31 (
// Equation(s):
// \pc_plus_4_D~31_combout  = (\pc_plus_4[30]~56_combout  & ((iwait) # (!\branch_or_jump~1_combout )))

	.dataa(gnd),
	.datab(iwait),
	.datac(\pc_plus_4[30]~56_combout ),
	.datad(\branch_or_jump~1_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_D~31_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_D~31 .lut_mask = 16'hC0F0;
defparam \pc_plus_4_D~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N5
dffeas \pc_plus_4_D[30] (
	.clk(CLK),
	.d(\pc_plus_4_D~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_D[30]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_D[30] .is_wysiwyg = "true";
defparam \pc_plus_4_D[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N12
cycloneive_lcell_comb \pc_plus_4_EX~31 (
// Equation(s):
// \pc_plus_4_EX~31_combout  = (\branch_or_jump~2_combout  & (pc_plus_4_D[30] & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\branch_or_jump~2_combout ),
	.datab(pc_plus_4_D[30]),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~31_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~31 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N13
dffeas \pc_plus_4_EX[30] (
	.clk(CLK),
	.d(\pc_plus_4_EX~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[30]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[30] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N4
cycloneive_lcell_comb \pc_plus_4_M~31 (
// Equation(s):
// \pc_plus_4_M~31_combout  = (pc_plus_4_EX[30] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_plus_4_EX[30]),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~31_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~31 .lut_mask = 16'h00F0;
defparam \pc_plus_4_M~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N5
dffeas \pc_plus_4_M[30] (
	.clk(CLK),
	.d(\pc_plus_4_M~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[30]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[30] .is_wysiwyg = "true";
defparam \pc_plus_4_M[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N2
cycloneive_lcell_comb \pc_plus_4_WB[30]~feeder (
// Equation(s):
// \pc_plus_4_WB[30]~feeder_combout  = pc_plus_4_M[30]

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pc_plus_4_M[30]),
	.cin(gnd),
	.combout(\pc_plus_4_WB[30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_WB[30]~feeder .lut_mask = 16'hFF00;
defparam \pc_plus_4_WB[30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N3
dffeas \pc_plus_4_WB[30] (
	.clk(CLK),
	.d(\pc_plus_4_WB[30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[30]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[30] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N20
cycloneive_lcell_comb \wdat_WB[30]~4 (
// Equation(s):
// \wdat_WB[30]~4_combout  = (\wdat_WB[28]~1_combout  & (\wdat_WB[28]~0_combout )) # (!\wdat_WB[28]~1_combout  & ((\wdat_WB[28]~0_combout  & ((pc_plus_4_WB[30]))) # (!\wdat_WB[28]~0_combout  & (porto_WB[30]))))

	.dataa(\wdat_WB[28]~1_combout ),
	.datab(\wdat_WB[28]~0_combout ),
	.datac(porto_WB[30]),
	.datad(pc_plus_4_WB[30]),
	.cin(gnd),
	.combout(\wdat_WB[30]~4_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[30]~4 .lut_mask = 16'hDC98;
defparam \wdat_WB[30]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N0
cycloneive_lcell_comb \wdat_WB[30]~5 (
// Equation(s):
// \wdat_WB[30]~5_combout  = (\wdat_WB[28]~1_combout  & ((\wdat_WB[30]~4_combout  & ((imm_WB[14]))) # (!\wdat_WB[30]~4_combout  & (dmemload_WB[30])))) # (!\wdat_WB[28]~1_combout  & (((\wdat_WB[30]~4_combout ))))

	.dataa(dmemload_WB[30]),
	.datab(imm_WB[14]),
	.datac(\wdat_WB[28]~1_combout ),
	.datad(\wdat_WB[30]~4_combout ),
	.cin(gnd),
	.combout(\wdat_WB[30]~5_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[30]~5 .lut_mask = 16'hCFA0;
defparam \wdat_WB[30]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N28
cycloneive_lcell_comb \sw_forwarding_output~1 (
// Equation(s):
// \sw_forwarding_output~1_combout  = (\lui_M~q  & ((imm_M[14]))) # (!\lui_M~q  & (porto_M_30))

	.dataa(gnd),
	.datab(porto_M_30),
	.datac(\lui_M~q ),
	.datad(imm_M[14]),
	.cin(gnd),
	.combout(\sw_forwarding_output~1_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~1 .lut_mask = 16'hFC0C;
defparam \sw_forwarding_output~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N18
cycloneive_lcell_comb \portB~18 (
// Equation(s):
// \portB~18_combout  = (\Equal3~2_combout  & (((\wdat_WB[30]~5_combout ) # (\portB~14_combout )))) # (!\Equal3~2_combout  & (rdata2_EX[30] & ((!\portB~14_combout ))))

	.dataa(rdata2_EX[30]),
	.datab(\wdat_WB[30]~5_combout ),
	.datac(\Equal3~2_combout ),
	.datad(\portB~14_combout ),
	.cin(gnd),
	.combout(\portB~18_combout ),
	.cout());
// synopsys translate_off
defparam \portB~18 .lut_mask = 16'hF0CA;
defparam \portB~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N6
cycloneive_lcell_comb \portB~19 (
// Equation(s):
// \portB~19_combout  = (\portB~14_combout  & ((\portB~18_combout  & (\sw_forwarding_output~1_combout )) # (!\portB~18_combout  & ((\sign_ext[16]~0_combout ))))) # (!\portB~14_combout  & (((\portB~18_combout ))))

	.dataa(\portB~14_combout ),
	.datab(\sw_forwarding_output~1_combout ),
	.datac(\sign_ext[16]~0_combout ),
	.datad(\portB~18_combout ),
	.cin(gnd),
	.combout(\portB~19_combout ),
	.cout());
// synopsys translate_off
defparam \portB~19 .lut_mask = 16'hDDA0;
defparam \portB~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N30
cycloneive_lcell_comb \portB~20 (
// Equation(s):
// \portB~20_combout  = (\portB~19_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q )))

	.dataa(\ShiftOp_EX~q ),
	.datab(\Equal3~2_combout ),
	.datac(gnd),
	.datad(\portB~19_combout ),
	.cin(gnd),
	.combout(\portB~20_combout ),
	.cout());
// synopsys translate_off
defparam \portB~20 .lut_mask = 16'hDD00;
defparam \portB~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N2
cycloneive_lcell_comb \rdata2_EX~2 (
// Equation(s):
// \rdata2_EX~2_combout  = (instruction_D[20] & (Mux33)) # (!instruction_D[20] & ((Mux331)))

	.dataa(instruction_D[20]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux33~9_combout ),
	.datad(\REGISTER_FILE|Mux33~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~2 .lut_mask = 16'hF5A0;
defparam \rdata2_EX~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N28
cycloneive_lcell_comb \rdata2_EX~3 (
// Equation(s):
// \rdata2_EX~3_combout  = (\always2~2_combout  & ((\rdata2_EX~2_combout ))) # (!\always2~2_combout  & (\portB~20_combout ))

	.dataa(gnd),
	.datab(\portB~20_combout ),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~2_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~3_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~3 .lut_mask = 16'hFC0C;
defparam \rdata2_EX~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N29
dffeas \rdata2_EX[30] (
	.clk(CLK),
	.d(\rdata2_EX~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[30]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[30] .is_wysiwyg = "true";
defparam \rdata2_EX[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N30
cycloneive_lcell_comb \rdata2_M~62 (
// Equation(s):
// \rdata2_M~62_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout )))) # (!\rdata2_M[16]~0_combout  & ((\rdata2_M[16]~1_combout  & ((\sw_forwarding_output~1_combout ))) # (!\rdata2_M[16]~1_combout  & (rdata2_EX[30]))))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(rdata2_EX[30]),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\sw_forwarding_output~1_combout ),
	.cin(gnd),
	.combout(\rdata2_M~62_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~62 .lut_mask = 16'hF4A4;
defparam \rdata2_M~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N22
cycloneive_lcell_comb \rdata2_M~63 (
// Equation(s):
// \rdata2_M~63_combout  = (\rdata2_M[16]~0_combout  & ((\rdata2_M~62_combout  & (\wdat_WB[30]~5_combout )) # (!\rdata2_M~62_combout  & ((ramiframload_30))))) # (!\rdata2_M[16]~0_combout  & (((\rdata2_M~62_combout ))))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(\wdat_WB[30]~5_combout ),
	.datac(\rdata2_M~62_combout ),
	.datad(\dpif.dmemload [30]),
	.cin(gnd),
	.combout(\rdata2_M~63_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~63 .lut_mask = 16'hDAD0;
defparam \rdata2_M~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N28
cycloneive_lcell_comb \imm_M~0 (
// Equation(s):
// \imm_M~0_combout  = (imm_EX[15] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(imm_EX[15]),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\imm_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \imm_M~0 .lut_mask = 16'h0C0C;
defparam \imm_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N29
dffeas \imm_M[15] (
	.clk(CLK),
	.d(\imm_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_M[15]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_M[15] .is_wysiwyg = "true";
defparam \imm_M[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N14
cycloneive_lcell_comb \imm_WB[15]~feeder (
// Equation(s):
// \imm_WB[15]~feeder_combout  = imm_M[15]

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(imm_M[15]),
	.cin(gnd),
	.combout(\imm_WB[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \imm_WB[15]~feeder .lut_mask = 16'hFF00;
defparam \imm_WB[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N15
dffeas \imm_WB[15] (
	.clk(CLK),
	.d(\imm_WB[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(imm_WB[15]),
	.prn(vcc));
// synopsys translate_off
defparam \imm_WB[15] .is_wysiwyg = "true";
defparam \imm_WB[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N18
cycloneive_lcell_comb \pc_plus_4_EX~30 (
// Equation(s):
// \pc_plus_4_EX~30_combout  = (pc_plus_4_D[31] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(pc_plus_4_D[31]),
	.datab(\branch_or_jump~2_combout ),
	.datac(\predicted_M~q ),
	.datad(\branch_taken~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_EX~30_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_EX~30 .lut_mask = 16'h8008;
defparam \pc_plus_4_EX~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N19
dffeas \pc_plus_4_EX[31] (
	.clk(CLK),
	.d(\pc_plus_4_EX~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_EX[31]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_EX[31] .is_wysiwyg = "true";
defparam \pc_plus_4_EX[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N26
cycloneive_lcell_comb \pc_plus_4_M~30 (
// Equation(s):
// \pc_plus_4_M~30_combout  = (pc_plus_4_EX[31] & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(pc_plus_4_EX[31]),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\pc_plus_4_M~30_combout ),
	.cout());
// synopsys translate_off
defparam \pc_plus_4_M~30 .lut_mask = 16'h00F0;
defparam \pc_plus_4_M~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N27
dffeas \pc_plus_4_M[31] (
	.clk(CLK),
	.d(\pc_plus_4_M~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_M[31]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_M[31] .is_wysiwyg = "true";
defparam \pc_plus_4_M[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N27
dffeas \pc_plus_4_WB[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(pc_plus_4_M[31]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_plus_4_WB[31]),
	.prn(vcc));
// synopsys translate_off
defparam \pc_plus_4_WB[31] .is_wysiwyg = "true";
defparam \pc_plus_4_WB[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N9
dffeas \dmemload_WB[31] (
	.clk(CLK),
	.d(\dpif.dmemload [31]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dmemload_WB[31]),
	.prn(vcc));
// synopsys translate_off
defparam \dmemload_WB[31] .is_wysiwyg = "true";
defparam \dmemload_WB[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N25
dffeas \porto_WB[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(porto_M_31),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(porto_WB[31]),
	.prn(vcc));
// synopsys translate_off
defparam \porto_WB[31] .is_wysiwyg = "true";
defparam \porto_WB[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N24
cycloneive_lcell_comb \wdat_WB[31]~2 (
// Equation(s):
// \wdat_WB[31]~2_combout  = (\wdat_WB[28]~1_combout  & ((dmemload_WB[31]) # ((\wdat_WB[28]~0_combout )))) # (!\wdat_WB[28]~1_combout  & (((porto_WB[31] & !\wdat_WB[28]~0_combout ))))

	.dataa(\wdat_WB[28]~1_combout ),
	.datab(dmemload_WB[31]),
	.datac(porto_WB[31]),
	.datad(\wdat_WB[28]~0_combout ),
	.cin(gnd),
	.combout(\wdat_WB[31]~2_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[31]~2 .lut_mask = 16'hAAD8;
defparam \wdat_WB[31]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N26
cycloneive_lcell_comb \wdat_WB[31]~3 (
// Equation(s):
// \wdat_WB[31]~3_combout  = (\wdat_WB[28]~0_combout  & ((\wdat_WB[31]~2_combout  & (imm_WB[15])) # (!\wdat_WB[31]~2_combout  & ((pc_plus_4_WB[31]))))) # (!\wdat_WB[28]~0_combout  & (((\wdat_WB[31]~2_combout ))))

	.dataa(\wdat_WB[28]~0_combout ),
	.datab(imm_WB[15]),
	.datac(pc_plus_4_WB[31]),
	.datad(\wdat_WB[31]~2_combout ),
	.cin(gnd),
	.combout(\wdat_WB[31]~3_combout ),
	.cout());
// synopsys translate_off
defparam \wdat_WB[31]~3 .lut_mask = 16'hDDA0;
defparam \wdat_WB[31]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N10
cycloneive_lcell_comb \sw_forwarding_output~0 (
// Equation(s):
// \sw_forwarding_output~0_combout  = (\lui_M~q  & (imm_M[15])) # (!\lui_M~q  & ((porto_M_31)))

	.dataa(gnd),
	.datab(imm_M[15]),
	.datac(\lui_M~q ),
	.datad(porto_M_31),
	.cin(gnd),
	.combout(\sw_forwarding_output~0_combout ),
	.cout());
// synopsys translate_off
defparam \sw_forwarding_output~0 .lut_mask = 16'hCFC0;
defparam \sw_forwarding_output~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N12
cycloneive_lcell_comb \rdata2_EX~0 (
// Equation(s):
// \rdata2_EX~0_combout  = (instruction_D[20] & (Mux32)) # (!instruction_D[20] & ((Mux321)))

	.dataa(gnd),
	.datab(\REGISTER_FILE|Mux32~9_combout ),
	.datac(instruction_D[20]),
	.datad(\REGISTER_FILE|Mux32~19_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~0 .lut_mask = 16'hCFC0;
defparam \rdata2_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N24
cycloneive_lcell_comb \rdata2_EX~1 (
// Equation(s):
// \rdata2_EX~1_combout  = (\always2~2_combout  & ((\rdata2_EX~0_combout ))) # (!\always2~2_combout  & (\portB~17_combout ))

	.dataa(\portB~17_combout ),
	.datab(gnd),
	.datac(\always2~2_combout ),
	.datad(\rdata2_EX~0_combout ),
	.cin(gnd),
	.combout(\rdata2_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_EX~1 .lut_mask = 16'hFA0A;
defparam \rdata2_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N25
dffeas \rdata2_EX[31] (
	.clk(CLK),
	.d(\rdata2_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata2_EX[31]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata2_EX[31] .is_wysiwyg = "true";
defparam \rdata2_EX[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N6
cycloneive_lcell_comb \rdata2_M~64 (
// Equation(s):
// \rdata2_M~64_combout  = (\rdata2_M[16]~0_combout  & (((\rdata2_M[16]~1_combout ) # (ramiframload_31)))) # (!\rdata2_M[16]~0_combout  & (rdata2_EX[31] & (!\rdata2_M[16]~1_combout )))

	.dataa(\rdata2_M[16]~0_combout ),
	.datab(rdata2_EX[31]),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\dpif.dmemload [31]),
	.cin(gnd),
	.combout(\rdata2_M~64_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~64 .lut_mask = 16'hAEA4;
defparam \rdata2_M~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N0
cycloneive_lcell_comb \rdata2_M~65 (
// Equation(s):
// \rdata2_M~65_combout  = (\rdata2_M[16]~1_combout  & ((\rdata2_M~64_combout  & (\wdat_WB[31]~3_combout )) # (!\rdata2_M~64_combout  & ((\sw_forwarding_output~0_combout ))))) # (!\rdata2_M[16]~1_combout  & (((\rdata2_M~64_combout ))))

	.dataa(\wdat_WB[31]~3_combout ),
	.datab(\sw_forwarding_output~0_combout ),
	.datac(\rdata2_M[16]~1_combout ),
	.datad(\rdata2_M~64_combout ),
	.cin(gnd),
	.combout(\rdata2_M~65_combout ),
	.cout());
// synopsys translate_off
defparam \rdata2_M~65 .lut_mask = 16'hAFC0;
defparam \rdata2_M~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N24
cycloneive_lcell_comb \porto_M~4 (
// Equation(s):
// \porto_M~4_combout  = (Selector30 & !\wsel_M~0_combout )

	.dataa(\ALU|Selector30~8_combout ),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\porto_M~4_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~4 .lut_mask = 16'h0A0A;
defparam \porto_M~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N0
cycloneive_lcell_comb \dWEN_M~0 (
// Equation(s):
// \dWEN_M~0_combout  = (\dWEN_EX~q  & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(\dWEN_EX~q ),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\dWEN_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \dWEN_M~0 .lut_mask = 16'h00CC;
defparam \dWEN_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N8
cycloneive_lcell_comb \dREN_EX~0 (
// Equation(s):
// \dREN_EX~0_combout  = (instruction_D[26] & (!instruction_D[30] & instruction_D[27])) # (!instruction_D[26] & (instruction_D[30] & !instruction_D[27]))

	.dataa(instruction_D[26]),
	.datab(instruction_D[30]),
	.datac(gnd),
	.datad(instruction_D[27]),
	.cin(gnd),
	.combout(\dREN_EX~0_combout ),
	.cout());
// synopsys translate_off
defparam \dREN_EX~0 .lut_mask = 16'h2244;
defparam \dREN_EX~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N16
cycloneive_lcell_comb \dREN_EX~1 (
// Equation(s):
// \dREN_EX~1_combout  = (instruction_D[31] & (\branch_or_jump~1_combout  & (\dREN_EX~0_combout  & Equal3)))

	.dataa(instruction_D[31]),
	.datab(\branch_or_jump~1_combout ),
	.datac(\dREN_EX~0_combout ),
	.datad(\CONTROL_UNIT|Equal3~1_combout ),
	.cin(gnd),
	.combout(\dREN_EX~1_combout ),
	.cout());
// synopsys translate_off
defparam \dREN_EX~1 .lut_mask = 16'h8000;
defparam \dREN_EX~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N17
dffeas dREN_EX(
	.clk(CLK),
	.d(\dREN_EX~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\dREN_EX~q ),
	.prn(vcc));
// synopsys translate_off
defparam dREN_EX.is_wysiwyg = "true";
defparam dREN_EX.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N30
cycloneive_lcell_comb \dREN_M~0 (
// Equation(s):
// \dREN_M~0_combout  = (\dREN_EX~q  & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\dREN_EX~q ),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\dREN_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \dREN_M~0 .lut_mask = 16'h00F0;
defparam \dREN_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N18
cycloneive_lcell_comb \instruction_D~76 (
// Equation(s):
// \instruction_D~76_combout  = (ramiframload_21 & (\branch_or_jump~1_combout  & iwait))

	.dataa(\dpif.dmemload [21]),
	.datab(\branch_or_jump~1_combout ),
	.datac(gnd),
	.datad(iwait),
	.cin(gnd),
	.combout(\instruction_D~76_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_D~76 .lut_mask = 16'h8800;
defparam \instruction_D~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N19
dffeas \instruction_D[21] (
	.clk(CLK),
	.d(\instruction_D~76_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_D[21]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_D[21] .is_wysiwyg = "true";
defparam \instruction_D[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N28
cycloneive_lcell_comb \instruction_EX~6 (
// Equation(s):
// \instruction_EX~6_combout  = (instruction_D[21] & (\branch_or_jump~2_combout  & (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(\predicted_M~q ),
	.datab(instruction_D[21]),
	.datac(\branch_taken~0_combout ),
	.datad(\branch_or_jump~2_combout ),
	.cin(gnd),
	.combout(\instruction_EX~6_combout ),
	.cout());
// synopsys translate_off
defparam \instruction_EX~6 .lut_mask = 16'h8400;
defparam \instruction_EX~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N29
dffeas \instruction_EX[21] (
	.clk(CLK),
	.d(\instruction_EX~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ALUSrc_EX~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instruction_EX[21]),
	.prn(vcc));
// synopsys translate_off
defparam \instruction_EX[21] .is_wysiwyg = "true";
defparam \instruction_EX[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N18
cycloneive_lcell_comb \rdata1_EX~64 (
// Equation(s):
// \rdata1_EX~64_combout  = (instruction_D[25] & ((Mux311))) # (!instruction_D[25] & (Mux312))

	.dataa(instruction_D[25]),
	.datab(gnd),
	.datac(\REGISTER_FILE|Mux31~19_combout ),
	.datad(\REGISTER_FILE|Mux31~9_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~64_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~64 .lut_mask = 16'hFA50;
defparam \rdata1_EX~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N16
cycloneive_lcell_comb \rdata1_EX~65 (
// Equation(s):
// \rdata1_EX~65_combout  = (\always2~2_combout  & ((\rdata1_EX~64_combout ))) # (!\always2~2_combout  & (\portA~69_combout ))

	.dataa(\portA~69_combout ),
	.datab(\always2~2_combout ),
	.datac(gnd),
	.datad(\rdata1_EX~64_combout ),
	.cin(gnd),
	.combout(\rdata1_EX~65_combout ),
	.cout());
// synopsys translate_off
defparam \rdata1_EX~65 .lut_mask = 16'hEE22;
defparam \rdata1_EX~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N17
dffeas \rdata1_EX[0] (
	.clk(CLK),
	.d(\rdata1_EX~65_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(!\branch_or_jump~1_combout ),
	.sload(gnd),
	.ena(\rdata1_EX[15]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(rdata1_EX[0]),
	.prn(vcc));
// synopsys translate_off
defparam \rdata1_EX[0] .is_wysiwyg = "true";
defparam \rdata1_EX[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N6
cycloneive_lcell_comb \regWrite_M~0 (
// Equation(s):
// \regWrite_M~0_combout  = (\RegWrite_EX~q  & !\wsel_M~0_combout )

	.dataa(\RegWrite_EX~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\regWrite_M~0_combout ),
	.cout());
// synopsys translate_off
defparam \regWrite_M~0 .lut_mask = 16'h00AA;
defparam \regWrite_M~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N7
dffeas regWrite_M(
	.clk(CLK),
	.d(\regWrite_M~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regWrite_M~q ),
	.prn(vcc));
// synopsys translate_off
defparam regWrite_M.is_wysiwyg = "true";
defparam regWrite_M.power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N21
dffeas regWrite_WB(
	.clk(CLK),
	.d(gnd),
	.asdata(\regWrite_M~q ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always4~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\regWrite_WB~q ),
	.prn(vcc));
// synopsys translate_off
defparam regWrite_WB.is_wysiwyg = "true";
defparam regWrite_WB.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N16
cycloneive_lcell_comb \portA~68 (
// Equation(s):
// \portA~68_combout  = (fuifforward_A_1 & ((\regWrite_WB~q  & (\wdat_WB[0]~61_combout )) # (!\regWrite_WB~q  & ((rdata1_EX[0]))))) # (!fuifforward_A_1 & (((rdata1_EX[0]))))

	.dataa(\wdat_WB[0]~61_combout ),
	.datab(rdata1_EX[0]),
	.datac(\FORWARDING_UNIT|fuif.forward_A[1]~5_combout ),
	.datad(\regWrite_WB~q ),
	.cin(gnd),
	.combout(\portA~68_combout ),
	.cout());
// synopsys translate_off
defparam \portA~68 .lut_mask = 16'hACCC;
defparam \portA~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N2
cycloneive_lcell_comb \portA~73 (
// Equation(s):
// \portA~73_combout  = (Equal3 & ((instruction_EX[21] & ((\portA~68_combout ))) # (!instruction_EX[21] & (rdata1_EX[0])))) # (!Equal3 & (((\portA~68_combout ))))

	.dataa(\FORWARDING_UNIT|Equal3~0_combout ),
	.datab(instruction_EX[21]),
	.datac(rdata1_EX[0]),
	.datad(\portA~68_combout ),
	.cin(gnd),
	.combout(\portA~73_combout ),
	.cout());
// synopsys translate_off
defparam \portA~73 .lut_mask = 16'hFD20;
defparam \portA~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N6
cycloneive_lcell_comb \portA~69 (
// Equation(s):
// \portA~69_combout  = (fuifforward_A_01 & (!\lui_M~q  & (porto_M_0))) # (!fuifforward_A_01 & (((\portA~73_combout ))))

	.dataa(\lui_M~q ),
	.datab(porto_M_0),
	.datac(\FORWARDING_UNIT|fuif.forward_A[0]~6_combout ),
	.datad(\portA~73_combout ),
	.cin(gnd),
	.combout(\portA~69_combout ),
	.cout());
// synopsys translate_off
defparam \portA~69 .lut_mask = 16'h4F40;
defparam \portA~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N14
cycloneive_lcell_comb \porto_M~35 (
// Equation(s):
// \porto_M~35_combout  = (Selector312) # ((!\portB~92_combout  & (!\portA~69_combout  & Selector0)))

	.dataa(\portB~92_combout ),
	.datab(\portA~69_combout ),
	.datac(\ALU|Selector31~8_combout ),
	.datad(\ALU|Selector0~5_combout ),
	.cin(gnd),
	.combout(\porto_M~35_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~35 .lut_mask = 16'hF1F0;
defparam \porto_M~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N0
cycloneive_lcell_comb \porto_M~5 (
// Equation(s):
// \porto_M~5_combout  = (!\wsel_M~0_combout  & ((Selector311) # ((\porto_M~35_combout ) # (Selector31))))

	.dataa(\ALU|Selector31~5_combout ),
	.datab(\wsel_M~0_combout ),
	.datac(\porto_M~35_combout ),
	.datad(\ALU|Selector31~4_combout ),
	.cin(gnd),
	.combout(\porto_M~5_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~5 .lut_mask = 16'h3332;
defparam \porto_M~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N8
cycloneive_lcell_comb \porto_M~6 (
// Equation(s):
// \porto_M~6_combout  = (!\wsel_M~0_combout  & Selector28)

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(\ALU|Selector28~10_combout ),
	.cin(gnd),
	.combout(\porto_M~6_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~6 .lut_mask = 16'h0F00;
defparam \porto_M~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N0
cycloneive_lcell_comb \porto_M~7 (
// Equation(s):
// \porto_M~7_combout  = (!\wsel_M~0_combout  & Selector29)

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(gnd),
	.datad(\ALU|Selector29~10_combout ),
	.cin(gnd),
	.combout(\porto_M~7_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~7 .lut_mask = 16'h3300;
defparam \porto_M~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N0
cycloneive_lcell_comb \porto_M~8 (
// Equation(s):
// \porto_M~8_combout  = (!\wsel_M~0_combout  & Selector26)

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(\ALU|Selector26~6_combout ),
	.cin(gnd),
	.combout(\porto_M~8_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~8 .lut_mask = 16'h0F00;
defparam \porto_M~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N0
cycloneive_lcell_comb \porto_M~36 (
// Equation(s):
// \porto_M~36_combout  = (!\wsel_M~0_combout  & ((Selector27) # ((Selector272) # (Selector271))))

	.dataa(\ALU|Selector27~0_combout ),
	.datab(\wsel_M~0_combout ),
	.datac(\ALU|Selector27~6_combout ),
	.datad(\ALU|Selector27~3_combout ),
	.cin(gnd),
	.combout(\porto_M~36_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~36 .lut_mask = 16'h3332;
defparam \porto_M~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N20
cycloneive_lcell_comb \porto_M~9 (
// Equation(s):
// \porto_M~9_combout  = (Selector24 & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ALU|Selector24~8_combout ),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\porto_M~9_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~9 .lut_mask = 16'h00F0;
defparam \porto_M~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N8
cycloneive_lcell_comb \porto_M~10 (
// Equation(s):
// \porto_M~10_combout  = (!\wsel_M~0_combout  & Selector25)

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(\ALU|Selector25~7_combout ),
	.cin(gnd),
	.combout(\porto_M~10_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~10 .lut_mask = 16'h0F00;
defparam \porto_M~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N12
cycloneive_lcell_comb \porto_M~11 (
// Equation(s):
// \porto_M~11_combout  = (!\wsel_M~0_combout  & Selector22)

	.dataa(\wsel_M~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ALU|Selector22~8_combout ),
	.cin(gnd),
	.combout(\porto_M~11_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~11 .lut_mask = 16'h5500;
defparam \porto_M~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N16
cycloneive_lcell_comb \porto_M~12 (
// Equation(s):
// \porto_M~12_combout  = (!\wsel_M~0_combout  & Selector23)

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(gnd),
	.datad(\ALU|Selector23~8_combout ),
	.cin(gnd),
	.combout(\porto_M~12_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~12 .lut_mask = 16'h3300;
defparam \porto_M~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N0
cycloneive_lcell_comb \porto_M~13 (
// Equation(s):
// \porto_M~13_combout  = (!\wsel_M~0_combout  & Selector20)

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(gnd),
	.datad(\ALU|Selector20~8_combout ),
	.cin(gnd),
	.combout(\porto_M~13_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~13 .lut_mask = 16'h3300;
defparam \porto_M~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N20
cycloneive_lcell_comb \porto_M~14 (
// Equation(s):
// \porto_M~14_combout  = (!\wsel_M~0_combout  & Selector21)

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(\ALU|Selector21~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\porto_M~14_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~14 .lut_mask = 16'h3030;
defparam \porto_M~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N18
cycloneive_lcell_comb \porto_M~15 (
// Equation(s):
// \porto_M~15_combout  = (!\wsel_M~0_combout  & Selector18)

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(\ALU|Selector18~7_combout ),
	.cin(gnd),
	.combout(\porto_M~15_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~15 .lut_mask = 16'h0F00;
defparam \porto_M~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N22
cycloneive_lcell_comb \porto_M~16 (
// Equation(s):
// \porto_M~16_combout  = (!\wsel_M~0_combout  & ((Selector19) # ((ShiftLeft0 & Selector16))))

	.dataa(\wsel_M~0_combout ),
	.datab(\ALU|ShiftLeft0~57_combout ),
	.datac(\ALU|Selector16~3_combout ),
	.datad(\ALU|Selector19~6_combout ),
	.cin(gnd),
	.combout(\porto_M~16_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~16 .lut_mask = 16'h5540;
defparam \porto_M~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N18
cycloneive_lcell_comb \porto_M~17 (
// Equation(s):
// \porto_M~17_combout  = (!\wsel_M~0_combout  & Selector161)

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(\ALU|Selector16~11_combout ),
	.cin(gnd),
	.combout(\porto_M~17_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~17 .lut_mask = 16'h0F00;
defparam \porto_M~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N28
cycloneive_lcell_comb \porto_M~18 (
// Equation(s):
// \porto_M~18_combout  = (Selector17 & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ALU|Selector17~8_combout ),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\porto_M~18_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~18 .lut_mask = 16'h00F0;
defparam \porto_M~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N10
cycloneive_lcell_comb \porto_M~19 (
// Equation(s):
// \porto_M~19_combout  = (!\wsel_M~0_combout  & Selector14)

	.dataa(\wsel_M~0_combout ),
	.datab(gnd),
	.datac(\ALU|Selector14~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\porto_M~19_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~19 .lut_mask = 16'h5050;
defparam \porto_M~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N20
cycloneive_lcell_comb \porto_M~20 (
// Equation(s):
// \porto_M~20_combout  = (!\wsel_M~0_combout  & Selector15)

	.dataa(\wsel_M~0_combout ),
	.datab(gnd),
	.datac(\ALU|Selector15~11_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\porto_M~20_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~20 .lut_mask = 16'h5050;
defparam \porto_M~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N16
cycloneive_lcell_comb \porto_M~21 (
// Equation(s):
// \porto_M~21_combout  = (Selector121 & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ALU|Selector12~18_combout ),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\porto_M~21_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~21 .lut_mask = 16'h00F0;
defparam \porto_M~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N18
cycloneive_lcell_comb \porto_M~22 (
// Equation(s):
// \porto_M~22_combout  = (Selector13 & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ALU|Selector13~8_combout ),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\porto_M~22_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~22 .lut_mask = 16'h00F0;
defparam \porto_M~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N6
cycloneive_lcell_comb \porto_M~23 (
// Equation(s):
// \porto_M~23_combout  = (Selector10 & !\wsel_M~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ALU|Selector10~8_combout ),
	.datad(\wsel_M~0_combout ),
	.cin(gnd),
	.combout(\porto_M~23_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~23 .lut_mask = 16'h00F0;
defparam \porto_M~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N14
cycloneive_lcell_comb \porto_M~24 (
// Equation(s):
// \porto_M~24_combout  = (!\wsel_M~0_combout  & Selector11)

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(gnd),
	.datad(\ALU|Selector11~8_combout ),
	.cin(gnd),
	.combout(\porto_M~24_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~24 .lut_mask = 16'h3300;
defparam \porto_M~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N28
cycloneive_lcell_comb \porto_M~25 (
// Equation(s):
// \porto_M~25_combout  = (!\wsel_M~0_combout  & ((Selector8) # ((Selector12 & ShiftRight0))))

	.dataa(\wsel_M~0_combout ),
	.datab(\ALU|Selector12~10_combout ),
	.datac(\ALU|ShiftRight0~91_combout ),
	.datad(\ALU|Selector8~7_combout ),
	.cin(gnd),
	.combout(\porto_M~25_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~25 .lut_mask = 16'h5540;
defparam \porto_M~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N14
cycloneive_lcell_comb \porto_M~26 (
// Equation(s):
// \porto_M~26_combout  = (!\wsel_M~0_combout  & Selector9)

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(\ALU|Selector9~8_combout ),
	.cin(gnd),
	.combout(\porto_M~26_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~26 .lut_mask = 16'h0F00;
defparam \porto_M~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N20
cycloneive_lcell_comb \porto_M~27 (
// Equation(s):
// \porto_M~27_combout  = (!\wsel_M~0_combout  & Selector62)

	.dataa(\wsel_M~0_combout ),
	.datab(gnd),
	.datac(\ALU|Selector6~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\porto_M~27_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~27 .lut_mask = 16'h5050;
defparam \porto_M~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N16
cycloneive_lcell_comb \porto_M~28 (
// Equation(s):
// \porto_M~28_combout  = (Selector7 & !\wsel_M~0_combout )

	.dataa(\ALU|Selector7~7_combout ),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\porto_M~28_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~28 .lut_mask = 16'h0A0A;
defparam \porto_M~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N18
cycloneive_lcell_comb \porto_M~29 (
// Equation(s):
// \porto_M~29_combout  = (!\wsel_M~0_combout  & Selector4)

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(\ALU|Selector4~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\porto_M~29_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~29 .lut_mask = 16'h3030;
defparam \porto_M~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N30
cycloneive_lcell_comb \porto_M~30 (
// Equation(s):
// \porto_M~30_combout  = (!\wsel_M~0_combout  & Selector5)

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(\ALU|Selector5~7_combout ),
	.cin(gnd),
	.combout(\porto_M~30_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~30 .lut_mask = 16'h0F00;
defparam \porto_M~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N16
cycloneive_lcell_comb \porto_M~31 (
// Equation(s):
// \porto_M~31_combout  = (!\wsel_M~0_combout  & Selector2)

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(gnd),
	.datad(\ALU|Selector2~11_combout ),
	.cin(gnd),
	.combout(\porto_M~31_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~31 .lut_mask = 16'h3300;
defparam \porto_M~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N14
cycloneive_lcell_comb \porto_M~32 (
// Equation(s):
// \porto_M~32_combout  = (!\wsel_M~0_combout  & Selector3)

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(gnd),
	.datad(\ALU|Selector3~9_combout ),
	.cin(gnd),
	.combout(\porto_M~32_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~32 .lut_mask = 16'h3300;
defparam \porto_M~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N30
cycloneive_lcell_comb \porto_M~33 (
// Equation(s):
// \porto_M~33_combout  = (!\wsel_M~0_combout  & Selector01)

	.dataa(gnd),
	.datab(gnd),
	.datac(\wsel_M~0_combout ),
	.datad(\ALU|Selector0~27_combout ),
	.cin(gnd),
	.combout(\porto_M~33_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~33 .lut_mask = 16'h0F00;
defparam \porto_M~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N2
cycloneive_lcell_comb \porto_M~34 (
// Equation(s):
// \porto_M~34_combout  = (!\wsel_M~0_combout  & Selector1)

	.dataa(gnd),
	.datab(\wsel_M~0_combout ),
	.datac(gnd),
	.datad(\ALU|Selector1~9_combout ),
	.cin(gnd),
	.combout(\porto_M~34_combout ),
	.cout());
// synopsys translate_off
defparam \porto_M~34 .lut_mask = 16'h3300;
defparam \porto_M~34 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module alu (
	ALUOp_EX_0,
	ALUOp_EX_1,
	ALUOp_EX_2,
	ALUOp_EX_3,
	ShiftOp_EX,
	portB,
	portB1,
	portB2,
	portB3,
	portB4,
	portB5,
	portB6,
	portB7,
	portB8,
	portB9,
	portB10,
	portB11,
	portB12,
	portB13,
	portB14,
	portB15,
	portB16,
	portB17,
	portB18,
	portB19,
	portB20,
	portB21,
	portB22,
	portB23,
	portB24,
	portB25,
	portB26,
	portB27,
	portB28,
	fuifforward_A_1,
	portA,
	portA1,
	portB29,
	portB30,
	portA2,
	wdat_WB_3,
	portA3,
	portA4,
	portB31,
	portA5,
	portA6,
	portA7,
	portA8,
	portB32,
	portA9,
	portA10,
	portA11,
	portA12,
	portA13,
	portA14,
	portA15,
	portA16,
	portB33,
	portA17,
	portA18,
	portA19,
	portA20,
	portA21,
	portA22,
	portA23,
	portA24,
	portA25,
	portA26,
	portA27,
	portA28,
	portA29,
	portA30,
	portA31,
	portA32,
	Selector0,
	Selector30,
	portB34,
	portB35,
	Selector31,
	Selector311,
	Selector312,
	Selector28,
	Selector29,
	Selector26,
	Selector27,
	Selector271,
	Selector272,
	Selector273,
	Selector24,
	Selector25,
	Selector22,
	Selector16,
	Selector23,
	Selector20,
	Selector21,
	Selector18,
	Selector19,
	ShiftLeft0,
	Selector161,
	Selector17,
	Selector12,
	Selector14,
	Selector15,
	Selector121,
	Selector13,
	Selector10,
	Selector11,
	Selector8,
	Selector9,
	Selector6,
	Selector61,
	Selector62,
	Selector7,
	Selector4,
	Selector5,
	Selector2,
	Selector3,
	Selector01,
	Selector1,
	Selector63,
	Selector64,
	Selector313,
	Equal3,
	ShiftRight0,
	devpor,
	devclrn,
	devoe);
input 	ALUOp_EX_0;
input 	ALUOp_EX_1;
input 	ALUOp_EX_2;
input 	ALUOp_EX_3;
input 	ShiftOp_EX;
input 	portB;
input 	portB1;
input 	portB2;
input 	portB3;
input 	portB4;
input 	portB5;
input 	portB6;
input 	portB7;
input 	portB8;
input 	portB9;
input 	portB10;
input 	portB11;
input 	portB12;
input 	portB13;
input 	portB14;
input 	portB15;
input 	portB16;
input 	portB17;
input 	portB18;
input 	portB19;
input 	portB20;
input 	portB21;
input 	portB22;
input 	portB23;
input 	portB24;
input 	portB25;
input 	portB26;
input 	portB27;
input 	portB28;
input 	fuifforward_A_1;
input 	portA;
input 	portA1;
input 	portB29;
input 	portB30;
input 	portA2;
input 	wdat_WB_3;
input 	portA3;
input 	portA4;
input 	portB31;
input 	portA5;
input 	portA6;
input 	portA7;
input 	portA8;
input 	portB32;
input 	portA9;
input 	portA10;
input 	portA11;
input 	portA12;
input 	portA13;
input 	portA14;
input 	portA15;
input 	portA16;
input 	portB33;
input 	portA17;
input 	portA18;
input 	portA19;
input 	portA20;
input 	portA21;
input 	portA22;
input 	portA23;
input 	portA24;
input 	portA25;
input 	portA26;
input 	portA27;
input 	portA28;
input 	portA29;
input 	portA30;
input 	portA31;
input 	portA32;
output 	Selector0;
output 	Selector30;
input 	portB34;
input 	portB35;
output 	Selector31;
output 	Selector311;
output 	Selector312;
output 	Selector28;
output 	Selector29;
output 	Selector26;
output 	Selector27;
output 	Selector271;
output 	Selector272;
output 	Selector273;
output 	Selector24;
output 	Selector25;
output 	Selector22;
output 	Selector16;
output 	Selector23;
output 	Selector20;
output 	Selector21;
output 	Selector18;
output 	Selector19;
output 	ShiftLeft0;
output 	Selector161;
output 	Selector17;
output 	Selector12;
output 	Selector14;
output 	Selector15;
output 	Selector121;
output 	Selector13;
output 	Selector10;
output 	Selector11;
output 	Selector8;
output 	Selector9;
output 	Selector6;
output 	Selector61;
output 	Selector62;
output 	Selector7;
output 	Selector4;
output 	Selector5;
output 	Selector2;
output 	Selector3;
output 	Selector01;
output 	Selector1;
output 	Selector63;
output 	Selector64;
output 	Selector313;
input 	Equal3;
output 	ShiftRight0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~12_combout ;
wire \Add1~16_combout ;
wire \ShiftLeft0~2_combout ;
wire \ShiftRight0~70_combout ;
wire \Selector29~1_combout ;
wire \ShiftLeft0~37_combout ;
wire \ShiftLeft0~46_combout ;
wire \ShiftLeft0~47_combout ;
wire \Selector21~3_combout ;
wire \Selector0~16_combout ;
wire \Selector8~2_combout ;
wire \Selector6~3_combout ;
wire \ShiftLeft0~91_combout ;
wire \ShiftLeft0~92_combout ;
wire \ShiftLeft0~94_combout ;
wire \Selector1~2_combout ;
wire \Selector1~3_combout ;
wire \Selector1~4_combout ;
wire \Selector0~4_combout ;
wire \Selector0~3_combout ;
wire \Selector30~3_combout ;
wire \Selector30~4_combout ;
wire \ShiftLeft0~13_combout ;
wire \ShiftLeft0~14_combout ;
wire \ShiftLeft0~4_combout ;
wire \ShiftLeft0~5_combout ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~6_combout ;
wire \ShiftLeft0~7_combout ;
wire \ShiftLeft0~9_combout ;
wire \ShiftLeft0~11_combout ;
wire \ShiftLeft0~12_combout ;
wire \Selector30~1_combout ;
wire \Selector30~2_combout ;
wire \Selector0~2_combout ;
wire \Selector30~5_combout ;
wire \Selector0~7_combout ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \Selector30~6_combout ;
wire \Selector30~7_combout ;
wire \Selector0~0_combout ;
wire \ShiftLeft0~8_combout ;
wire \ShiftLeft0~10_combout ;
wire \Selector31~0_combout ;
wire \ShiftRight0~13_combout ;
wire \ShiftRight0~12_combout ;
wire \ShiftRight0~14_combout ;
wire \ShiftRight0~15_combout ;
wire \ShiftRight0~6_combout ;
wire \ShiftRight0~5_combout ;
wire \ShiftRight0~7_combout ;
wire \ShiftRight0~3_combout ;
wire \ShiftRight0~2_combout ;
wire \ShiftRight0~4_combout ;
wire \ShiftRight0~8_combout ;
wire \ShiftRight0~16_combout ;
wire \ShiftRight0~20_combout ;
wire \ShiftRight0~19_combout ;
wire \ShiftRight0~21_combout ;
wire \ShiftRight0~17_combout ;
wire \ShiftRight0~18_combout ;
wire \ShiftRight0~22_combout ;
wire \ShiftRight0~26_combout ;
wire \ShiftRight0~27_combout ;
wire \ShiftRight0~28_combout ;
wire \ShiftRight0~24_combout ;
wire \ShiftRight0~23_combout ;
wire \ShiftRight0~25_combout ;
wire \Selector22~0_combout ;
wire \ShiftRight0~29_combout ;
wire \Selector30~0_combout ;
wire \Add0~0_combout ;
wire \Selector0~6_combout ;
wire \Add1~0_combout ;
wire \Selector31~2_combout ;
wire \Selector31~3_combout ;
wire \LessThan1~1_cout ;
wire \LessThan1~3_cout ;
wire \LessThan1~5_cout ;
wire \LessThan1~7_cout ;
wire \LessThan1~9_cout ;
wire \LessThan1~11_cout ;
wire \LessThan1~13_cout ;
wire \LessThan1~15_cout ;
wire \LessThan1~17_cout ;
wire \LessThan1~19_cout ;
wire \LessThan1~21_cout ;
wire \LessThan1~23_cout ;
wire \LessThan1~25_cout ;
wire \LessThan1~27_cout ;
wire \LessThan1~29_cout ;
wire \LessThan1~31_cout ;
wire \LessThan1~33_cout ;
wire \LessThan1~35_cout ;
wire \LessThan1~37_cout ;
wire \LessThan1~39_cout ;
wire \LessThan1~41_cout ;
wire \LessThan1~43_cout ;
wire \LessThan1~45_cout ;
wire \LessThan1~47_cout ;
wire \LessThan1~49_cout ;
wire \LessThan1~51_cout ;
wire \LessThan1~53_cout ;
wire \LessThan1~55_cout ;
wire \LessThan1~57_cout ;
wire \LessThan1~59_cout ;
wire \LessThan1~61_cout ;
wire \LessThan1~62_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~23_cout ;
wire \LessThan0~25_cout ;
wire \LessThan0~27_cout ;
wire \LessThan0~29_cout ;
wire \LessThan0~31_cout ;
wire \LessThan0~33_cout ;
wire \LessThan0~35_cout ;
wire \LessThan0~37_cout ;
wire \LessThan0~39_cout ;
wire \LessThan0~41_cout ;
wire \LessThan0~43_cout ;
wire \LessThan0~45_cout ;
wire \LessThan0~47_cout ;
wire \LessThan0~49_cout ;
wire \LessThan0~51_cout ;
wire \LessThan0~53_cout ;
wire \LessThan0~55_cout ;
wire \LessThan0~57_cout ;
wire \LessThan0~59_cout ;
wire \LessThan0~61_cout ;
wire \LessThan0~62_combout ;
wire \Selector31~1_combout ;
wire \ShiftRight0~40_combout ;
wire \ShiftRight0~41_combout ;
wire \ShiftRight0~42_combout ;
wire \ShiftRight0~38_combout ;
wire \ShiftRight0~37_combout ;
wire \ShiftRight0~39_combout ;
wire \ShiftRight0~43_combout ;
wire \ShiftRight0~31_combout ;
wire \ShiftRight0~30_combout ;
wire \ShiftRight0~32_combout ;
wire \ShiftRight0~36_combout ;
wire \ShiftRight0~44_combout ;
wire \ShiftRight0~53_combout ;
wire \ShiftRight0~52_combout ;
wire \ShiftRight0~54_combout ;
wire \Selector23~0_combout ;
wire \ShiftRight0~48_combout ;
wire \ShiftRight0~49_combout ;
wire \ShiftRight0~50_combout ;
wire \ShiftRight0~46_combout ;
wire \ShiftRight0~45_combout ;
wire \ShiftRight0~47_combout ;
wire \ShiftRight0~51_combout ;
wire \ShiftRight0~58_combout ;
wire \ShiftLeft0~15_combout ;
wire \Selector31~7_combout ;
wire \Selector0~10_combout ;
wire \Selector0~8_combout ;
wire \Selector28~4_combout ;
wire \Selector28~5_combout ;
wire \ShiftLeft0~17_combout ;
wire \ShiftLeft0~16_combout ;
wire \Selector29~0_combout ;
wire \ShiftLeft0~18_combout ;
wire \ShiftLeft0~19_combout ;
wire \Selector0~13_combout ;
wire \Selector28~7_combout ;
wire \Selector0~11_combout ;
wire \Add0~3 ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~6_combout ;
wire \Selector28~6_combout ;
wire \Selector28~8_combout ;
wire \Selector28~9_combout ;
wire \Selector12~4_combout ;
wire \Selector12~5_combout ;
wire \Selector16~0_combout ;
wire \ShiftRight0~67_combout ;
wire \ShiftRight0~68_combout ;
wire \Selector20~0_combout ;
wire \ShiftRight0~63_combout ;
wire \ShiftRight0~64_combout ;
wire \ShiftRight0~65_combout ;
wire \ShiftRight0~66_combout ;
wire \ShiftRight0~69_combout ;
wire \Selector12~19_combout ;
wire \Selector28~0_combout ;
wire \ShiftRight0~59_combout ;
wire \Selector2~2_combout ;
wire \Selector28~1_combout ;
wire \ShiftRight0~9_combout ;
wire \ShiftRight0~60_combout ;
wire \ShiftRight0~10_combout ;
wire \ShiftRight0~61_combout ;
wire \ShiftRight0~62_combout ;
wire \Selector28~2_combout ;
wire \Selector28~3_combout ;
wire \ShiftRight0~34_combout ;
wire \ShiftRight0~72_combout ;
wire \ShiftRight0~71_combout ;
wire \ShiftRight0~73_combout ;
wire \Selector29~2_combout ;
wire \Selector29~3_combout ;
wire \ShiftRight0~74_combout ;
wire \ShiftRight0~75_combout ;
wire \ShiftRight0~76_combout ;
wire \ShiftRight0~55_combout ;
wire \ShiftRight0~77_combout ;
wire \Selector21~0_combout ;
wire \ShiftRight0~78_combout ;
wire \ShiftLeft0~20_combout ;
wire \ShiftLeft0~21_combout ;
wire \Selector0~9_combout ;
wire \Selector29~4_combout ;
wire \Selector29~5_combout ;
wire \Selector29~6_combout ;
wire \Add1~4_combout ;
wire \Add0~4_combout ;
wire \Selector29~7_combout ;
wire \Selector29~8_combout ;
wire \Selector29~9_combout ;
wire \Selector26~2_combout ;
wire \Selector26~0_combout ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \Add0~7 ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \Selector26~1_combout ;
wire \Selector0~1_combout ;
wire \Selector24~0_combout ;
wire \ShiftLeft0~22_combout ;
wire \ShiftLeft0~23_combout ;
wire \ShiftLeft0~24_combout ;
wire \Selector4~0_combout ;
wire \ShiftRight0~80_combout ;
wire \ShiftRight0~81_combout ;
wire \ShiftRight0~11_combout ;
wire \ShiftRight0~79_combout ;
wire \Selector26~3_combout ;
wire \Selector26~4_combout ;
wire \Selector26~5_combout ;
wire \Add0~8_combout ;
wire \Add1~8_combout ;
wire \ShiftLeft0~25_combout ;
wire \ShiftLeft0~27_combout ;
wire \ShiftLeft0~26_combout ;
wire \ShiftLeft0~28_combout ;
wire \ShiftLeft0~29_combout ;
wire \Selector4~1_combout ;
wire \ShiftRight0~56_combout ;
wire \ShiftRight0~57_combout ;
wire \ShiftRight0~82_combout ;
wire \ShiftRight0~33_combout ;
wire \ShiftRight0~35_combout ;
wire \Selector27~1_combout ;
wire \ShiftRight0~83_combout ;
wire \ShiftRight0~84_combout ;
wire \Selector27~2_combout ;
wire \Selector27~4_combout ;
wire \Selector27~5_combout ;
wire \ShiftRight0~85_combout ;
wire \Selector24~6_combout ;
wire \Selector24~7_combout ;
wire \Selector24~1_combout ;
wire \Selector24~3_combout ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~14_combout ;
wire \Add0~11 ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \Selector24~2_combout ;
wire \Selector24~4_combout ;
wire \ShiftLeft0~30_combout ;
wire \ShiftLeft0~31_combout ;
wire \ShiftLeft0~32_combout ;
wire \Selector4~2_combout ;
wire \Selector24~5_combout ;
wire \Selector25~2_combout ;
wire \Selector25~0_combout ;
wire \Add0~12_combout ;
wire \Selector25~1_combout ;
wire \Selector25~3_combout ;
wire \ShiftRight0~89_combout ;
wire \Selector4~3_combout ;
wire \ShiftRight0~88_combout ;
wire \ShiftRight0~90_combout ;
wire \ShiftRight0~87_combout ;
wire \Selector25~5_combout ;
wire \Selector25~6_combout ;
wire \ShiftLeft0~35_combout ;
wire \Selector25~4_combout ;
wire \Selector0~12_combout ;
wire \Add0~15 ;
wire \Add0~17 ;
wire \Add0~18_combout ;
wire \Selector22~7_combout ;
wire \ShiftLeft0~38_combout ;
wire \ShiftLeft0~39_combout ;
wire \ShiftLeft0~36_combout ;
wire \ShiftLeft0~40_combout ;
wire \Selector22~5_combout ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~18_combout ;
wire \Selector22~6_combout ;
wire \Selector22~3_combout ;
wire \Selector22~2_combout ;
wire \Selector16~1_combout ;
wire \Selector16~2_combout ;
wire \Selector22~4_combout ;
wire \Selector20~1_combout ;
wire \Selector12~6_combout ;
wire \Selector22~1_combout ;
wire \Selector0~14_combout ;
wire \ShiftLeft0~41_combout ;
wire \ShiftLeft0~42_combout ;
wire \ShiftLeft0~33_combout ;
wire \ShiftLeft0~43_combout ;
wire \Selector23~1_combout ;
wire \Add0~16_combout ;
wire \Selector23~3_combout ;
wire \Selector23~2_combout ;
wire \Selector23~4_combout ;
wire \Selector23~5_combout ;
wire \Selector23~6_combout ;
wire \Selector23~7_combout ;
wire \Add0~19 ;
wire \Add0~21 ;
wire \Add0~22_combout ;
wire \Selector20~2_combout ;
wire \Selector20~3_combout ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~22_combout ;
wire \Selector20~4_combout ;
wire \Selector20~5_combout ;
wire \Selector20~6_combout ;
wire \Selector20~7_combout ;
wire \Add0~20_combout ;
wire \Selector21~4_combout ;
wire \ShiftLeft0~34_combout ;
wire \ShiftLeft0~48_combout ;
wire \ShiftLeft0~49_combout ;
wire \ShiftLeft0~50_combout ;
wire \ShiftLeft0~51_combout ;
wire \Selector21~5_combout ;
wire \Add1~20_combout ;
wire \Selector21~2_combout ;
wire \Selector21~6_combout ;
wire \Selector21~1_combout ;
wire \Selector18~0_combout ;
wire \Selector18~2_combout ;
wire \Selector18~3_combout ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~26_combout ;
wire \Selector18~4_combout ;
wire \ShiftLeft0~52_combout ;
wire \ShiftLeft0~44_combout ;
wire \ShiftLeft0~53_combout ;
wire \Selector10~0_combout ;
wire \ShiftLeft0~54_combout ;
wire \Selector18~1_combout ;
wire \Add0~23 ;
wire \Add0~25 ;
wire \Add0~26_combout ;
wire \Selector18~5_combout ;
wire \Selector18~6_combout ;
wire \Add0~24_combout ;
wire \Selector19~3_combout ;
wire \Selector19~4_combout ;
wire \Add1~24_combout ;
wire \Selector19~5_combout ;
wire \Selector19~0_combout ;
wire \Selector19~1_combout ;
wire \Selector19~2_combout ;
wire \ShiftLeft0~55_combout ;
wire \ShiftLeft0~56_combout ;
wire \Selector11~0_combout ;
wire \Add0~27 ;
wire \Add0~29 ;
wire \Add0~30_combout ;
wire \Selector16~4_combout ;
wire \Selector16~5_combout ;
wire \Selector16~6_combout ;
wire \ShiftLeft0~58_combout ;
wire \ShiftLeft0~59_combout ;
wire \ShiftLeft0~45_combout ;
wire \Selector8~0_combout ;
wire \ShiftLeft0~60_combout ;
wire \Selector16~7_combout ;
wire \Selector16~8_combout ;
wire \Selector16~9_combout ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~30_combout ;
wire \Selector16~10_combout ;
wire \Selector17~9_combout ;
wire \ShiftLeft0~61_combout ;
wire \ShiftLeft0~62_combout ;
wire \Selector9~0_combout ;
wire \ShiftLeft0~63_combout ;
wire \Selector17~2_combout ;
wire \Selector17~4_combout ;
wire \Add1~28_combout ;
wire \Selector17~3_combout ;
wire \Selector17~5_combout ;
wire \Add0~28_combout ;
wire \Selector17~6_combout ;
wire \Selector17~7_combout ;
wire \Selector0~15_combout ;
wire \Add0~31 ;
wire \Add0~33 ;
wire \Add0~34_combout ;
wire \Selector14~1_combout ;
wire \Selector14~0_combout ;
wire \Selector12~7_combout ;
wire \Selector14~2_combout ;
wire \ShiftLeft0~64_combout ;
wire \ShiftLeft0~65_combout ;
wire \ShiftLeft0~66_combout ;
wire \Selector12~8_combout ;
wire \Selector12~9_combout ;
wire \Selector14~3_combout ;
wire \Selector14~4_combout ;
wire \Selector12~11_combout ;
wire \Selector14~5_combout ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~34_combout ;
wire \Selector14~6_combout ;
wire \Selector15~9_combout ;
wire \Add1~32_combout ;
wire \Selector15~10_combout ;
wire \Add0~32_combout ;
wire \Selector15~5_combout ;
wire \Selector15~4_combout ;
wire \Selector15~6_combout ;
wire \ShiftLeft0~67_combout ;
wire \ShiftLeft0~68_combout ;
wire \Selector15~12_combout ;
wire \Selector15~7_combout ;
wire \Selector15~8_combout ;
wire \Selector12~20_combout ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~38_combout ;
wire \Selector12~17_combout ;
wire \Add0~35 ;
wire \Add0~37 ;
wire \Add0~38_combout ;
wire \Selector12~12_combout ;
wire \Selector12~13_combout ;
wire \Selector12~14_combout ;
wire \ShiftLeft0~70_combout ;
wire \ShiftLeft0~71_combout ;
wire \ShiftLeft0~72_combout ;
wire \Selector12~15_combout ;
wire \Selector12~16_combout ;
wire \Add0~36_combout ;
wire \Selector13~2_combout ;
wire \Selector13~3_combout ;
wire \Selector13~4_combout ;
wire \Selector13~9_combout ;
wire \Selector13~5_combout ;
wire \Add1~36_combout ;
wire \Selector13~6_combout ;
wire \Selector13~7_combout ;
wire \Add0~39 ;
wire \Add0~41 ;
wire \Add0~42_combout ;
wire \Selector10~1_combout ;
wire \Selector10~2_combout ;
wire \Selector10~3_combout ;
wire \Selector10~4_combout ;
wire \Selector10~5_combout ;
wire \Selector10~6_combout ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~42_combout ;
wire \Selector10~7_combout ;
wire \Add0~40_combout ;
wire \Selector11~2_combout ;
wire \Selector11~1_combout ;
wire \Selector11~4_combout ;
wire \Selector11~3_combout ;
wire \Selector11~5_combout ;
wire \Add1~40_combout ;
wire \Selector11~6_combout ;
wire \Selector11~7_combout ;
wire \Selector8~1_combout ;
wire \Selector8~5_combout ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~46_combout ;
wire \Selector8~3_combout ;
wire \Selector8~4_combout ;
wire \Selector8~6_combout ;
wire \Add0~43 ;
wire \Add0~45 ;
wire \Add0~46_combout ;
wire \Add0~44_combout ;
wire \ShiftLeft0~85_combout ;
wire \ShiftLeft0~80_combout ;
wire \ShiftLeft0~86_combout ;
wire \ShiftLeft0~74_combout ;
wire \Selector1~0_combout ;
wire \Selector9~6_combout ;
wire \Add1~44_combout ;
wire \Selector9~7_combout ;
wire \Selector9~1_combout ;
wire \Selector9~2_combout ;
wire \Selector9~3_combout ;
wire \Selector9~4_combout ;
wire \Selector9~5_combout ;
wire \Add0~47 ;
wire \Add0~49 ;
wire \Add0~50_combout ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~50_combout ;
wire \Selector4~4_combout ;
wire \ShiftLeft0~83_combout ;
wire \ShiftLeft0~87_combout ;
wire \ShiftLeft0~88_combout ;
wire \ShiftLeft0~76_combout ;
wire \ShiftLeft0~77_combout ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \Selector6~4_combout ;
wire \Selector6~6_combout ;
wire \Add0~48_combout ;
wire \Selector7~0_combout ;
wire \Selector7~1_combout ;
wire \ShiftLeft0~79_combout ;
wire \ShiftLeft0~81_combout ;
wire \ShiftLeft0~69_combout ;
wire \ShiftLeft0~89_combout ;
wire \ShiftLeft0~90_combout ;
wire \Selector7~2_combout ;
wire \ShiftLeft0~97_combout ;
wire \Selector7~3_combout ;
wire \Selector7~4_combout ;
wire \Selector7~5_combout ;
wire \Add1~48_combout ;
wire \Selector7~6_combout ;
wire \Add0~51 ;
wire \Add0~53 ;
wire \Add0~54_combout ;
wire \Selector4~10_combout ;
wire \Add1~51 ;
wire \Add1~53 ;
wire \Add1~54_combout ;
wire \Selector4~11_combout ;
wire \Selector4~5_combout ;
wire \Selector4~8_combout ;
wire \ShiftLeft0~84_combout ;
wire \Selector4~6_combout ;
wire \Selector4~7_combout ;
wire \Selector4~9_combout ;
wire \Selector5~0_combout ;
wire \Selector5~1_combout ;
wire \ShiftLeft0~73_combout ;
wire \ShiftLeft0~75_combout ;
wire \Selector5~2_combout ;
wire \Selector5~3_combout ;
wire \Selector5~4_combout ;
wire \Add0~52_combout ;
wire \Selector5~5_combout ;
wire \Add1~52_combout ;
wire \Selector5~6_combout ;
wire \Add0~55 ;
wire \Add0~57 ;
wire \Add0~58_combout ;
wire \Selector2~3_combout ;
wire \Selector2~9_combout ;
wire \ShiftLeft0~78_combout ;
wire \Selector2~4_combout ;
wire \Selector2~5_combout ;
wire \Selector2~6_combout ;
wire \Selector2~7_combout ;
wire \Selector2~12_combout ;
wire \Selector2~8_combout ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~58_combout ;
wire \Selector2~10_combout ;
wire \Selector3~2_combout ;
wire \Add0~56_combout ;
wire \Selector3~7_combout ;
wire \Selector3~10_combout ;
wire \ShiftLeft0~93_combout ;
wire \ShiftLeft0~96_combout ;
wire \Selector3~3_combout ;
wire \ShiftLeft0~82_combout ;
wire \Selector3~4_combout ;
wire \Selector3~5_combout ;
wire \Selector3~6_combout ;
wire \Add1~56_combout ;
wire \Selector3~8_combout ;
wire \Add0~59 ;
wire \Add0~61 ;
wire \Add0~62_combout ;
wire \Selector0~17_combout ;
wire \Selector0~18_combout ;
wire \Selector0~19_combout ;
wire \Add1~59 ;
wire \Add1~61 ;
wire \Add1~62_combout ;
wire \Selector0~20_combout ;
wire \Selector0~21_combout ;
wire \ShiftLeft0~95_combout ;
wire \Selector0~22_combout ;
wire \Selector0~23_combout ;
wire \Selector0~24_combout ;
wire \Selector0~25_combout ;
wire \Selector0~26_combout ;
wire \Selector1~1_combout ;
wire \Add0~60_combout ;
wire \Selector1~7_combout ;
wire \Selector1~5_combout ;
wire \Selector1~6_combout ;
wire \Add1~60_combout ;
wire \Selector1~8_combout ;
wire \Selector7~8_combout ;
wire \Selector31~6_combout ;
wire \ShiftRight0~86_combout ;


// Location: LCCOMB_X58_Y31_N12
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((\portB~84_combout  $ (\portA~21_combout  $ (\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((\portB~84_combout  & (\portA~21_combout  & !\Add1~11 )) # (!\portB~84_combout  & ((\portA~21_combout ) # (!\Add1~11 ))))

	.dataa(portB27),
	.datab(portA7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h964D;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N16
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((\portB~76_combout  $ (\portA~17_combout  $ (\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((\portB~76_combout  & (\portA~17_combout  & !\Add1~15 )) # (!\portB~76_combout  & ((\portA~17_combout ) # (!\Add1~15 ))))

	.dataa(portB23),
	.datab(portA5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h964D;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N26
cycloneive_lcell_comb \ShiftLeft0~2 (
// Equation(s):
// \ShiftLeft0~2_combout  = (\portB~20_combout ) # ((\portB~23_combout ) # ((\portB~17_combout ) # (\portB~26_combout )))

	.dataa(portB1),
	.datab(portB2),
	.datac(portB),
	.datad(portB3),
	.cin(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~2 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N8
cycloneive_lcell_comb \ShiftRight0~70 (
// Equation(s):
// \ShiftRight0~70_combout  = (\portB~97_combout  & ((\ShiftRight0~41_combout ))) # (!\portB~97_combout  & (\ShiftRight0~33_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftRight0~33_combout ),
	.datad(\ShiftRight0~41_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~70 .lut_mask = 16'hFA50;
defparam \ShiftRight0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N10
cycloneive_lcell_comb \Selector29~1 (
// Equation(s):
// \Selector29~1_combout  = (\Selector2~2_combout  & (((!\ShiftLeft0~17_combout )))) # (!\Selector2~2_combout  & ((\ShiftLeft0~17_combout  & (\ShiftRight0~31_combout )) # (!\ShiftLeft0~17_combout  & ((\ShiftRight0~70_combout )))))

	.dataa(\Selector2~2_combout ),
	.datab(\ShiftRight0~31_combout ),
	.datac(\ShiftRight0~70_combout ),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\Selector29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~1 .lut_mask = 16'h44FA;
defparam \Selector29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N10
cycloneive_lcell_comb \ShiftLeft0~37 (
// Equation(s):
// \ShiftLeft0~37_combout  = (!\portB~97_combout  & (!\portB~100_combout  & (\ShiftLeft0~13_combout  & \portB~103_combout )))

	.dataa(portB30),
	.datab(portB31),
	.datac(\ShiftLeft0~13_combout ),
	.datad(portB32),
	.cin(gnd),
	.combout(\ShiftLeft0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~37 .lut_mask = 16'h1000;
defparam \ShiftLeft0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N12
cycloneive_lcell_comb \ShiftLeft0~46 (
// Equation(s):
// \ShiftLeft0~46_combout  = (!\portB~103_combout  & ((\portB~100_combout  & (\ShiftLeft0~31_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~45_combout )))))

	.dataa(portB31),
	.datab(portB32),
	.datac(\ShiftLeft0~31_combout ),
	.datad(\ShiftLeft0~45_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~46 .lut_mask = 16'h3120;
defparam \ShiftLeft0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N26
cycloneive_lcell_comb \ShiftLeft0~47 (
// Equation(s):
// \ShiftLeft0~47_combout  = (\ShiftLeft0~46_combout ) # ((!\portB~100_combout  & (\portB~103_combout  & \ShiftLeft0~19_combout )))

	.dataa(portB31),
	.datab(portB32),
	.datac(\ShiftLeft0~19_combout ),
	.datad(\ShiftLeft0~46_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~47 .lut_mask = 16'hFF40;
defparam \ShiftLeft0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N16
cycloneive_lcell_comb \Selector21~3 (
// Equation(s):
// \Selector21~3_combout  = (\portA~36_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \portB~109_combout )))) # (!\portA~36_combout  & (((\Selector0~8_combout  & \portB~109_combout ))))

	.dataa(\Selector0~9_combout ),
	.datab(portA15),
	.datac(\Selector0~8_combout ),
	.datad(portB35),
	.cin(gnd),
	.combout(\Selector21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~3 .lut_mask = 16'hF8C0;
defparam \Selector21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N12
cycloneive_lcell_comb \Selector0~16 (
// Equation(s):
// \Selector0~16_combout  = (\portB~100_combout  & (\ShiftLeft0~71_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~84_combout )))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftLeft0~71_combout ),
	.datad(\ShiftLeft0~84_combout ),
	.cin(gnd),
	.combout(\Selector0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~16 .lut_mask = 16'hF3C0;
defparam \Selector0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N30
cycloneive_lcell_comb \Selector8~2 (
// Equation(s):
// \Selector8~2_combout  = (\Selector12~5_combout  & (!\Selector12~8_combout  & \Selector0~16_combout ))

	.dataa(gnd),
	.datab(\Selector12~5_combout ),
	.datac(\Selector12~8_combout ),
	.datad(\Selector0~16_combout ),
	.cin(gnd),
	.combout(\Selector8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~2 .lut_mask = 16'h0C00;
defparam \Selector8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N26
cycloneive_lcell_comb \Selector6~3 (
// Equation(s):
// \Selector6~3_combout  = (!\portB~107_combout  & (\ShiftRight0~22_combout  & (!\portB~103_combout  & !\ShiftLeft0~16_combout )))

	.dataa(portB33),
	.datab(\ShiftRight0~22_combout ),
	.datac(portB32),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~3 .lut_mask = 16'h0004;
defparam \Selector6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N30
cycloneive_lcell_comb \ShiftLeft0~91 (
// Equation(s):
// \ShiftLeft0~91_combout  = (\portB~92_combout  & ((\portA~49_combout ))) # (!\portB~92_combout  & (\portA~47_combout ))

	.dataa(gnd),
	.datab(portA21),
	.datac(portA22),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~91 .lut_mask = 16'hF0CC;
defparam \ShiftLeft0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N16
cycloneive_lcell_comb \ShiftLeft0~92 (
// Equation(s):
// \ShiftLeft0~92_combout  = (\portB~97_combout  & ((\ShiftLeft0~87_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~91_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftLeft0~91_combout ),
	.datad(\ShiftLeft0~87_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~92 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N18
cycloneive_lcell_comb \ShiftLeft0~94 (
// Equation(s):
// \ShiftLeft0~94_combout  = (\portB~97_combout  & (\ShiftLeft0~89_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~93_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~89_combout ),
	.datac(portB30),
	.datad(\ShiftLeft0~93_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~94 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N14
cycloneive_lcell_comb \Selector1~2 (
// Equation(s):
// \Selector1~2_combout  = (\portA~43_combout  & (((\Selector0~10_combout  & !\portB~20_combout )))) # (!\portA~43_combout  & ((\portB~20_combout  & ((\Selector0~10_combout ))) # (!\portB~20_combout  & (\Selector0~13_combout ))))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~10_combout ),
	.datac(portA19),
	.datad(portB1),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~2 .lut_mask = 16'h0CCA;
defparam \Selector1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N20
cycloneive_lcell_comb \Selector1~3 (
// Equation(s):
// \Selector1~3_combout  = (\ShiftLeft0~14_combout  & (((\Selector0~21_combout ) # (\ShiftLeft0~96_combout )))) # (!\ShiftLeft0~14_combout  & (\portA~43_combout  & (!\Selector0~21_combout )))

	.dataa(portA19),
	.datab(\ShiftLeft0~14_combout ),
	.datac(\Selector0~21_combout ),
	.datad(\ShiftLeft0~96_combout ),
	.cin(gnd),
	.combout(\Selector1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~3 .lut_mask = 16'hCEC2;
defparam \Selector1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N6
cycloneive_lcell_comb \Selector1~4 (
// Equation(s):
// \Selector1~4_combout  = (\Selector0~21_combout  & ((\Selector1~3_combout  & (\ShiftLeft0~94_combout )) # (!\Selector1~3_combout  & ((\portA~41_combout ))))) # (!\Selector0~21_combout  & (((\Selector1~3_combout ))))

	.dataa(\ShiftLeft0~94_combout ),
	.datab(portA18),
	.datac(\Selector0~21_combout ),
	.datad(\Selector1~3_combout ),
	.cin(gnd),
	.combout(\Selector1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~4 .lut_mask = 16'hAFC0;
defparam \Selector1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N6
cycloneive_lcell_comb \Selector0~5 (
// Equation(s):
// Selector0 = (ALUOp_EX[0] & (ALUOp_EX[2] & (!ALUOp_EX[3] & ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(Selector0),
	.cout());
// synopsys translate_off
defparam \Selector0~5 .lut_mask = 16'h0800;
defparam \Selector0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N30
cycloneive_lcell_comb \Selector30~8 (
// Equation(s):
// Selector30 = (\Selector30~4_combout ) # ((\Selector30~2_combout ) # ((\Selector30~7_combout ) # (\Selector30~0_combout )))

	.dataa(\Selector30~4_combout ),
	.datab(\Selector30~2_combout ),
	.datac(\Selector30~7_combout ),
	.datad(\Selector30~0_combout ),
	.cin(gnd),
	.combout(Selector30),
	.cout());
// synopsys translate_off
defparam \Selector30~8 .lut_mask = 16'hFFFE;
defparam \Selector30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N20
cycloneive_lcell_comb \Selector31~4 (
// Equation(s):
// Selector31 = (\Selector31~3_combout ) # ((ALUOp_EX[3] & (!ALUOp_EX[2] & \Selector31~1_combout )))

	.dataa(ALUOp_EX_3),
	.datab(ALUOp_EX_2),
	.datac(\Selector31~3_combout ),
	.datad(\Selector31~1_combout ),
	.cin(gnd),
	.combout(Selector31),
	.cout());
// synopsys translate_off
defparam \Selector31~4 .lut_mask = 16'hF2F0;
defparam \Selector31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N10
cycloneive_lcell_comb \Selector31~5 (
// Equation(s):
// Selector311 = (\Selector31~0_combout  & ((\ShiftRight0~44_combout ) # ((\portB~107_combout  & \ShiftRight0~58_combout ))))

	.dataa(portB33),
	.datab(\Selector31~0_combout ),
	.datac(\ShiftRight0~44_combout ),
	.datad(\ShiftRight0~58_combout ),
	.cin(gnd),
	.combout(Selector311),
	.cout());
// synopsys translate_off
defparam \Selector31~5 .lut_mask = 16'hC8C0;
defparam \Selector31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N8
cycloneive_lcell_comb \Selector31~8 (
// Equation(s):
// Selector312 = (\portA~69_combout  & ((\Selector31~7_combout ) # ((!\ShiftLeft0~15_combout  & \Selector30~1_combout ))))

	.dataa(\ShiftLeft0~15_combout ),
	.datab(\Selector31~7_combout ),
	.datac(portA32),
	.datad(\Selector30~1_combout ),
	.cin(gnd),
	.combout(Selector312),
	.cout());
// synopsys translate_off
defparam \Selector31~8 .lut_mask = 16'hD0C0;
defparam \Selector31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N0
cycloneive_lcell_comb \Selector28~10 (
// Equation(s):
// Selector28 = (\Selector28~9_combout ) # ((\Selector28~3_combout ) # ((\Selector16~0_combout  & \ShiftRight0~69_combout )))

	.dataa(\Selector28~9_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\ShiftRight0~69_combout ),
	.datad(\Selector28~3_combout ),
	.cin(gnd),
	.combout(Selector28),
	.cout());
// synopsys translate_off
defparam \Selector28~10 .lut_mask = 16'hFFEA;
defparam \Selector28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N16
cycloneive_lcell_comb \Selector29~10 (
// Equation(s):
// Selector29 = (\Selector29~3_combout ) # ((\Selector29~9_combout ) # ((\Selector16~0_combout  & \ShiftRight0~78_combout )))

	.dataa(\Selector16~0_combout ),
	.datab(\Selector29~3_combout ),
	.datac(\ShiftRight0~78_combout ),
	.datad(\Selector29~9_combout ),
	.cin(gnd),
	.combout(Selector29),
	.cout());
// synopsys translate_off
defparam \Selector29~10 .lut_mask = 16'hFFEC;
defparam \Selector29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N20
cycloneive_lcell_comb \Selector26~6 (
// Equation(s):
// Selector26 = (\Selector26~2_combout ) # ((\Selector26~0_combout ) # ((\Selector26~1_combout ) # (\Selector26~5_combout )))

	.dataa(\Selector26~2_combout ),
	.datab(\Selector26~0_combout ),
	.datac(\Selector26~1_combout ),
	.datad(\Selector26~5_combout ),
	.cin(gnd),
	.combout(Selector26),
	.cout());
// synopsys translate_off
defparam \Selector26~6 .lut_mask = 16'hFFFE;
defparam \Selector26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N8
cycloneive_lcell_comb \Selector27~0 (
// Equation(s):
// Selector27 = (\Selector0~7_combout  & ((\Add0~8_combout ) # ((\Selector0~6_combout  & \Add1~8_combout )))) # (!\Selector0~7_combout  & (\Selector0~6_combout  & ((\Add1~8_combout ))))

	.dataa(\Selector0~7_combout ),
	.datab(\Selector0~6_combout ),
	.datac(\Add0~8_combout ),
	.datad(\Add1~8_combout ),
	.cin(gnd),
	.combout(Selector27),
	.cout());
// synopsys translate_off
defparam \Selector27~0 .lut_mask = 16'hECA0;
defparam \Selector27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N10
cycloneive_lcell_comb \Selector27~3 (
// Equation(s):
// Selector271 = (\Selector31~0_combout  & ((\Selector27~2_combout ) # ((\Selector24~0_combout  & \ShiftLeft0~29_combout )))) # (!\Selector31~0_combout  & (\Selector24~0_combout  & (\ShiftLeft0~29_combout )))

	.dataa(\Selector31~0_combout ),
	.datab(\Selector24~0_combout ),
	.datac(\ShiftLeft0~29_combout ),
	.datad(\Selector27~2_combout ),
	.cin(gnd),
	.combout(Selector271),
	.cout());
// synopsys translate_off
defparam \Selector27~3 .lut_mask = 16'hEAC0;
defparam \Selector27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N30
cycloneive_lcell_comb \Selector27~6 (
// Equation(s):
// Selector272 = (\Selector27~5_combout  & ((\Selector0~4_combout ) # ((\Selector0~2_combout )))) # (!\Selector27~5_combout  & (((\Selector27~4_combout ))))

	.dataa(\Selector0~4_combout ),
	.datab(\Selector27~4_combout ),
	.datac(\Selector0~2_combout ),
	.datad(\Selector27~5_combout ),
	.cin(gnd),
	.combout(Selector272),
	.cout());
// synopsys translate_off
defparam \Selector27~6 .lut_mask = 16'hFACC;
defparam \Selector27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N8
cycloneive_lcell_comb \Selector27~7 (
// Equation(s):
// Selector273 = (Selector272) # ((Selector27) # (Selector271))

	.dataa(gnd),
	.datab(Selector272),
	.datac(Selector27),
	.datad(Selector271),
	.cin(gnd),
	.combout(Selector273),
	.cout());
// synopsys translate_off
defparam \Selector27~7 .lut_mask = 16'hFFFC;
defparam \Selector27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N16
cycloneive_lcell_comb \Selector24~8 (
// Equation(s):
// Selector24 = (\Selector24~4_combout ) # ((\Selector24~5_combout ) # ((\Selector24~7_combout  & \Selector31~0_combout )))

	.dataa(\Selector24~7_combout ),
	.datab(\Selector31~0_combout ),
	.datac(\Selector24~4_combout ),
	.datad(\Selector24~5_combout ),
	.cin(gnd),
	.combout(Selector24),
	.cout());
// synopsys translate_off
defparam \Selector24~8 .lut_mask = 16'hFFF8;
defparam \Selector24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N6
cycloneive_lcell_comb \Selector25~7 (
// Equation(s):
// Selector25 = (\Selector25~3_combout ) # ((\Selector25~4_combout ) # ((\Selector25~6_combout  & \Selector31~0_combout )))

	.dataa(\Selector25~3_combout ),
	.datab(\Selector25~6_combout ),
	.datac(\Selector31~0_combout ),
	.datad(\Selector25~4_combout ),
	.cin(gnd),
	.combout(Selector25),
	.cout());
// synopsys translate_off
defparam \Selector25~7 .lut_mask = 16'hFFEA;
defparam \Selector25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N16
cycloneive_lcell_comb \Selector22~8 (
// Equation(s):
// Selector22 = (\Selector22~7_combout ) # ((\Selector22~6_combout ) # ((\Selector22~4_combout ) # (\Selector22~1_combout )))

	.dataa(\Selector22~7_combout ),
	.datab(\Selector22~6_combout ),
	.datac(\Selector22~4_combout ),
	.datad(\Selector22~1_combout ),
	.cin(gnd),
	.combout(Selector22),
	.cout());
// synopsys translate_off
defparam \Selector22~8 .lut_mask = 16'hFFFE;
defparam \Selector22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N20
cycloneive_lcell_comb \Selector16~3 (
// Equation(s):
// Selector16 = (\Selector0~14_combout  & (!\portB~107_combout  & (!\ShiftLeft0~12_combout  & !\ShiftLeft0~6_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(portB33),
	.datac(\ShiftLeft0~12_combout ),
	.datad(\ShiftLeft0~6_combout ),
	.cin(gnd),
	.combout(Selector16),
	.cout());
// synopsys translate_off
defparam \Selector16~3 .lut_mask = 16'h0002;
defparam \Selector16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N24
cycloneive_lcell_comb \Selector23~8 (
// Equation(s):
// Selector23 = (\Selector23~1_combout ) # ((\Selector23~7_combout ) # ((\Selector20~1_combout  & \ShiftRight0~51_combout )))

	.dataa(\Selector20~1_combout ),
	.datab(\ShiftRight0~51_combout ),
	.datac(\Selector23~1_combout ),
	.datad(\Selector23~7_combout ),
	.cin(gnd),
	.combout(Selector23),
	.cout());
// synopsys translate_off
defparam \Selector23~8 .lut_mask = 16'hFFF8;
defparam \Selector23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N6
cycloneive_lcell_comb \Selector20~8 (
// Equation(s):
// Selector20 = (\Selector20~4_combout ) # ((\Selector20~7_combout ) # ((\Add0~22_combout  & \Selector0~12_combout )))

	.dataa(\Add0~22_combout ),
	.datab(\Selector20~4_combout ),
	.datac(\Selector0~12_combout ),
	.datad(\Selector20~7_combout ),
	.cin(gnd),
	.combout(Selector20),
	.cout());
// synopsys translate_off
defparam \Selector20~8 .lut_mask = 16'hFFEC;
defparam \Selector20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N4
cycloneive_lcell_comb \Selector21~7 (
// Equation(s):
// Selector21 = (\Selector21~6_combout ) # ((\Selector21~1_combout ) # ((\Add0~20_combout  & \Selector0~12_combout )))

	.dataa(\Add0~20_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Selector21~6_combout ),
	.datad(\Selector21~1_combout ),
	.cin(gnd),
	.combout(Selector21),
	.cout());
// synopsys translate_off
defparam \Selector21~7 .lut_mask = 16'hFFF8;
defparam \Selector21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N6
cycloneive_lcell_comb \Selector18~7 (
// Equation(s):
// Selector18 = (\Selector18~0_combout ) # ((\Selector18~4_combout ) # ((\Selector18~1_combout ) # (\Selector18~6_combout )))

	.dataa(\Selector18~0_combout ),
	.datab(\Selector18~4_combout ),
	.datac(\Selector18~1_combout ),
	.datad(\Selector18~6_combout ),
	.cin(gnd),
	.combout(Selector18),
	.cout());
// synopsys translate_off
defparam \Selector18~7 .lut_mask = 16'hFFFE;
defparam \Selector18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N16
cycloneive_lcell_comb \Selector19~6 (
// Equation(s):
// Selector19 = (\Selector19~5_combout ) # ((\Selector19~2_combout ) # ((\Selector0~12_combout  & \Add0~24_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Add0~24_combout ),
	.datac(\Selector19~5_combout ),
	.datad(\Selector19~2_combout ),
	.cin(gnd),
	.combout(Selector19),
	.cout());
// synopsys translate_off
defparam \Selector19~6 .lut_mask = 16'hFFF8;
defparam \Selector19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N10
cycloneive_lcell_comb \ShiftLeft0~57 (
// Equation(s):
// ShiftLeft0 = (\portB~103_combout  & (\ShiftLeft0~29_combout )) # (!\portB~103_combout  & ((\Selector11~0_combout )))

	.dataa(portB32),
	.datab(gnd),
	.datac(\ShiftLeft0~29_combout ),
	.datad(\Selector11~0_combout ),
	.cin(gnd),
	.combout(ShiftLeft0),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~57 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N20
cycloneive_lcell_comb \Selector16~11 (
// Equation(s):
// Selector161 = (\Selector16~8_combout ) # ((\Selector16~10_combout ) # ((\Add0~30_combout  & \Selector0~12_combout )))

	.dataa(\Add0~30_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Selector16~8_combout ),
	.datad(\Selector16~10_combout ),
	.cin(gnd),
	.combout(Selector161),
	.cout());
// synopsys translate_off
defparam \Selector16~11 .lut_mask = 16'hFFF8;
defparam \Selector16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N14
cycloneive_lcell_comb \Selector17~8 (
// Equation(s):
// Selector17 = (\Selector17~9_combout ) # ((\Selector17~2_combout ) # ((\Selector17~5_combout ) # (\Selector17~7_combout )))

	.dataa(\Selector17~9_combout ),
	.datab(\Selector17~2_combout ),
	.datac(\Selector17~5_combout ),
	.datad(\Selector17~7_combout ),
	.cin(gnd),
	.combout(Selector17),
	.cout());
// synopsys translate_off
defparam \Selector17~8 .lut_mask = 16'hFFFE;
defparam \Selector17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N0
cycloneive_lcell_comb \Selector12~10 (
// Equation(s):
// Selector12 = (\Selector0~15_combout  & (!\ShiftLeft0~12_combout  & (!\portB~107_combout  & !\ShiftLeft0~6_combout )))

	.dataa(\Selector0~15_combout ),
	.datab(\ShiftLeft0~12_combout ),
	.datac(portB33),
	.datad(\ShiftLeft0~6_combout ),
	.cin(gnd),
	.combout(Selector12),
	.cout());
// synopsys translate_off
defparam \Selector12~10 .lut_mask = 16'h0002;
defparam \Selector12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N28
cycloneive_lcell_comb \Selector14~7 (
// Equation(s):
// Selector14 = (\Selector14~4_combout ) # ((\Selector14~6_combout ) # ((\Add0~34_combout  & \Selector0~12_combout )))

	.dataa(\Add0~34_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Selector14~4_combout ),
	.datad(\Selector14~6_combout ),
	.cin(gnd),
	.combout(Selector14),
	.cout());
// synopsys translate_off
defparam \Selector14~7 .lut_mask = 16'hFFF8;
defparam \Selector14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N22
cycloneive_lcell_comb \Selector15~11 (
// Equation(s):
// Selector15 = (\Selector15~10_combout ) # ((\Selector15~8_combout ) # ((\Selector0~12_combout  & \Add0~32_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector15~10_combout ),
	.datac(\Add0~32_combout ),
	.datad(\Selector15~8_combout ),
	.cin(gnd),
	.combout(Selector15),
	.cout());
// synopsys translate_off
defparam \Selector15~11 .lut_mask = 16'hFFEC;
defparam \Selector15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N26
cycloneive_lcell_comb \Selector12~18 (
// Equation(s):
// Selector121 = (\Selector12~17_combout ) # ((\Selector12~16_combout ) # ((\Selector0~12_combout  & \Add0~38_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector12~17_combout ),
	.datac(\Add0~38_combout ),
	.datad(\Selector12~16_combout ),
	.cin(gnd),
	.combout(Selector121),
	.cout());
// synopsys translate_off
defparam \Selector12~18 .lut_mask = 16'hFFEC;
defparam \Selector12~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N20
cycloneive_lcell_comb \Selector13~8 (
// Equation(s):
// Selector13 = (\Selector13~5_combout ) # ((\Selector13~7_combout ) # ((\Selector0~12_combout  & \Add0~36_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Add0~36_combout ),
	.datac(\Selector13~5_combout ),
	.datad(\Selector13~7_combout ),
	.cin(gnd),
	.combout(Selector13),
	.cout());
// synopsys translate_off
defparam \Selector13~8 .lut_mask = 16'hFFF8;
defparam \Selector13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N4
cycloneive_lcell_comb \Selector10~8 (
// Equation(s):
// Selector10 = (\Selector10~5_combout ) # ((\Selector10~7_combout ) # ((\Add0~42_combout  & \Selector0~12_combout )))

	.dataa(\Add0~42_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Selector10~5_combout ),
	.datad(\Selector10~7_combout ),
	.cin(gnd),
	.combout(Selector10),
	.cout());
// synopsys translate_off
defparam \Selector10~8 .lut_mask = 16'hFFF8;
defparam \Selector10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N18
cycloneive_lcell_comb \Selector11~8 (
// Equation(s):
// Selector11 = (\Selector11~5_combout ) # ((\Selector11~7_combout ) # ((\Selector0~12_combout  & \Add0~40_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Add0~40_combout ),
	.datac(\Selector11~5_combout ),
	.datad(\Selector11~7_combout ),
	.cin(gnd),
	.combout(Selector11),
	.cout());
// synopsys translate_off
defparam \Selector11~8 .lut_mask = 16'hFFF8;
defparam \Selector11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N4
cycloneive_lcell_comb \Selector8~7 (
// Equation(s):
// Selector8 = (\Selector8~1_combout ) # ((\Selector8~6_combout ) # ((\Selector0~12_combout  & \Add0~46_combout )))

	.dataa(\Selector8~1_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Selector8~6_combout ),
	.datad(\Add0~46_combout ),
	.cin(gnd),
	.combout(Selector8),
	.cout());
// synopsys translate_off
defparam \Selector8~7 .lut_mask = 16'hFEFA;
defparam \Selector8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N24
cycloneive_lcell_comb \Selector9~8 (
// Equation(s):
// Selector9 = (\Selector9~7_combout ) # ((\Selector9~5_combout ) # ((\Selector0~12_combout  & \Add0~44_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Add0~44_combout ),
	.datac(\Selector9~7_combout ),
	.datad(\Selector9~5_combout ),
	.cin(gnd),
	.combout(Selector9),
	.cout());
// synopsys translate_off
defparam \Selector9~8 .lut_mask = 16'hFFF8;
defparam \Selector9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N14
cycloneive_lcell_comb \Selector6~0 (
// Equation(s):
// Selector6 = (\portB~35_combout  & ((\Selector0~2_combout ) # ((\Selector0~3_combout  & \portA~51_combout )))) # (!\portB~35_combout  & (((\portA~51_combout  & \Selector0~2_combout ))))

	.dataa(\Selector0~3_combout ),
	.datab(portB6),
	.datac(portA23),
	.datad(\Selector0~2_combout ),
	.cin(gnd),
	.combout(Selector6),
	.cout());
// synopsys translate_off
defparam \Selector6~0 .lut_mask = 16'hFC80;
defparam \Selector6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N14
cycloneive_lcell_comb \Selector6~5 (
// Equation(s):
// Selector61 = (\portA~51_combout  & (((\Selector0~4_combout  & !\portB~35_combout )))) # (!\portA~51_combout  & ((\portB~35_combout  & ((\Selector0~4_combout ))) # (!\portB~35_combout  & (Selector0))))

	.dataa(Selector0),
	.datab(\Selector0~4_combout ),
	.datac(portA23),
	.datad(portB6),
	.cin(gnd),
	.combout(Selector61),
	.cout());
// synopsys translate_off
defparam \Selector6~5 .lut_mask = 16'h0CCA;
defparam \Selector6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N24
cycloneive_lcell_comb \Selector6~7 (
// Equation(s):
// Selector62 = (Selector6) # ((\Selector6~6_combout ) # ((\Selector0~7_combout  & \Add0~50_combout )))

	.dataa(\Selector0~7_combout ),
	.datab(Selector6),
	.datac(\Add0~50_combout ),
	.datad(\Selector6~6_combout ),
	.cin(gnd),
	.combout(Selector62),
	.cout());
// synopsys translate_off
defparam \Selector6~7 .lut_mask = 16'hFFEC;
defparam \Selector6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N26
cycloneive_lcell_comb \Selector7~7 (
// Equation(s):
// Selector7 = (\Selector7~4_combout ) # ((\Selector7~6_combout ) # ((\Selector0~7_combout  & \Add0~48_combout )))

	.dataa(\Selector0~7_combout ),
	.datab(\Add0~48_combout ),
	.datac(\Selector7~4_combout ),
	.datad(\Selector7~6_combout ),
	.cin(gnd),
	.combout(Selector7),
	.cout());
// synopsys translate_off
defparam \Selector7~7 .lut_mask = 16'hFFF8;
defparam \Selector7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N8
cycloneive_lcell_comb \Selector4~12 (
// Equation(s):
// Selector4 = (\Selector4~11_combout ) # ((\Selector4~9_combout ) # ((\Selector0~7_combout  & \Add0~54_combout )))

	.dataa(\Selector0~7_combout ),
	.datab(\Add0~54_combout ),
	.datac(\Selector4~11_combout ),
	.datad(\Selector4~9_combout ),
	.cin(gnd),
	.combout(Selector4),
	.cout());
// synopsys translate_off
defparam \Selector4~12 .lut_mask = 16'hFFF8;
defparam \Selector4~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N10
cycloneive_lcell_comb \Selector5~7 (
// Equation(s):
// Selector5 = (\Selector5~4_combout ) # ((\Selector5~6_combout ) # ((\Selector0~7_combout  & \Add0~52_combout )))

	.dataa(\Selector0~7_combout ),
	.datab(\Selector5~4_combout ),
	.datac(\Add0~52_combout ),
	.datad(\Selector5~6_combout ),
	.cin(gnd),
	.combout(Selector5),
	.cout());
// synopsys translate_off
defparam \Selector5~7 .lut_mask = 16'hFFEC;
defparam \Selector5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N16
cycloneive_lcell_comb \Selector2~11 (
// Equation(s):
// Selector2 = (\Selector2~3_combout ) # ((\Selector2~10_combout ) # ((\Selector0~12_combout  & \Add0~58_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Add0~58_combout ),
	.datac(\Selector2~3_combout ),
	.datad(\Selector2~10_combout ),
	.cin(gnd),
	.combout(Selector2),
	.cout());
// synopsys translate_off
defparam \Selector2~11 .lut_mask = 16'hFFF8;
defparam \Selector2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N24
cycloneive_lcell_comb \Selector3~9 (
// Equation(s):
// Selector3 = (\Selector3~2_combout ) # ((\Selector3~8_combout ) # ((\Selector0~12_combout  & \Add0~56_combout )))

	.dataa(\Selector3~2_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Add0~56_combout ),
	.datad(\Selector3~8_combout ),
	.cin(gnd),
	.combout(Selector3),
	.cout());
// synopsys translate_off
defparam \Selector3~9 .lut_mask = 16'hFFEA;
defparam \Selector3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N16
cycloneive_lcell_comb \Selector0~27 (
// Equation(s):
// Selector01 = (\Selector0~17_combout ) # ((\Selector0~26_combout ) # ((\Selector0~12_combout  & \Add0~62_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Add0~62_combout ),
	.datac(\Selector0~17_combout ),
	.datad(\Selector0~26_combout ),
	.cin(gnd),
	.combout(Selector01),
	.cout());
// synopsys translate_off
defparam \Selector0~27 .lut_mask = 16'hFFF8;
defparam \Selector0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N10
cycloneive_lcell_comb \Selector1~9 (
// Equation(s):
// Selector1 = (\Selector1~1_combout ) # ((\Selector1~8_combout ) # ((\Selector0~12_combout  & \Add0~60_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector1~1_combout ),
	.datac(\Add0~60_combout ),
	.datad(\Selector1~8_combout ),
	.cin(gnd),
	.combout(Selector1),
	.cout());
// synopsys translate_off
defparam \Selector1~9 .lut_mask = 16'hFFEC;
defparam \Selector1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N22
cycloneive_lcell_comb \Selector6~8 (
// Equation(s):
// Selector63 = (\Add1~50_combout  & ((\Selector0~6_combout ) # ((\Selector0~7_combout  & \Add0~50_combout )))) # (!\Add1~50_combout  & (((\Selector0~7_combout  & \Add0~50_combout ))))

	.dataa(\Add1~50_combout ),
	.datab(\Selector0~6_combout ),
	.datac(\Selector0~7_combout ),
	.datad(\Add0~50_combout ),
	.cin(gnd),
	.combout(Selector63),
	.cout());
// synopsys translate_off
defparam \Selector6~8 .lut_mask = 16'hF888;
defparam \Selector6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N20
cycloneive_lcell_comb \Selector6~9 (
// Equation(s):
// Selector64 = (\Selector7~8_combout  & ((\ShiftRight0~22_combout ) # ((\Selector4~4_combout  & \Selector6~2_combout )))) # (!\Selector7~8_combout  & (\Selector4~4_combout  & ((\Selector6~2_combout ))))

	.dataa(\Selector7~8_combout ),
	.datab(\Selector4~4_combout ),
	.datac(\ShiftRight0~22_combout ),
	.datad(\Selector6~2_combout ),
	.cin(gnd),
	.combout(Selector64),
	.cout());
// synopsys translate_off
defparam \Selector6~9 .lut_mask = 16'hECA0;
defparam \Selector6~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N28
cycloneive_lcell_comb \Selector31~9 (
// Equation(s):
// Selector313 = (Selector311) # ((\Selector31~6_combout ) # ((Selector312) # (Selector31)))

	.dataa(Selector311),
	.datab(\Selector31~6_combout ),
	.datac(Selector312),
	.datad(Selector31),
	.cin(gnd),
	.combout(Selector313),
	.cout());
// synopsys translate_off
defparam \Selector31~9 .lut_mask = 16'hFFFE;
defparam \Selector31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N30
cycloneive_lcell_comb \ShiftRight0~91 (
// Equation(s):
// ShiftRight0 = (\ShiftRight0~86_combout ) # ((!\portB~100_combout  & (\ShiftRight0~67_combout  & !\portB~103_combout )))

	.dataa(portB31),
	.datab(\ShiftRight0~67_combout ),
	.datac(portB32),
	.datad(\ShiftRight0~86_combout ),
	.cin(gnd),
	.combout(ShiftRight0),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~91 .lut_mask = 16'hFF04;
defparam \ShiftRight0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N20
cycloneive_lcell_comb \Selector0~4 (
// Equation(s):
// \Selector0~4_combout  = (!ALUOp_EX[0] & (ALUOp_EX[2] & (!ALUOp_EX[3] & ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~4 .lut_mask = 16'h0400;
defparam \Selector0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N12
cycloneive_lcell_comb \Selector0~3 (
// Equation(s):
// \Selector0~3_combout  = (!ALUOp_EX[3] & (ALUOp_EX[2] & (!ALUOp_EX[0] & !ALUOp_EX[1])))

	.dataa(ALUOp_EX_3),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_0),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~3 .lut_mask = 16'h0004;
defparam \Selector0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N4
cycloneive_lcell_comb \Selector30~3 (
// Equation(s):
// \Selector30~3_combout  = (\portA~12_combout  & ((\Selector0~2_combout ) # ((\Selector0~3_combout  & \portB~97_combout ))))

	.dataa(\Selector0~2_combout ),
	.datab(\Selector0~3_combout ),
	.datac(portA1),
	.datad(portB30),
	.cin(gnd),
	.combout(\Selector30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~3 .lut_mask = 16'hE0A0;
defparam \Selector30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N12
cycloneive_lcell_comb \Selector30~4 (
// Equation(s):
// \Selector30~4_combout  = (\Selector30~3_combout ) # ((\Selector0~4_combout  & (\portA~12_combout  $ (\portB~97_combout ))))

	.dataa(\Selector0~4_combout ),
	.datab(portA1),
	.datac(portB30),
	.datad(\Selector30~3_combout ),
	.cin(gnd),
	.combout(\Selector30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~4 .lut_mask = 16'hFF28;
defparam \Selector30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N14
cycloneive_lcell_comb \ShiftLeft0~13 (
// Equation(s):
// \ShiftLeft0~13_combout  = (\portB~92_combout  & (\portA~69_combout )) # (!\portB~92_combout  & ((\portA~12_combout )))

	.dataa(portA32),
	.datab(gnd),
	.datac(portB29),
	.datad(portA1),
	.cin(gnd),
	.combout(\ShiftLeft0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~13 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N16
cycloneive_lcell_comb \ShiftLeft0~14 (
// Equation(s):
// \ShiftLeft0~14_combout  = (\portB~97_combout ) # (\portB~100_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(portB30),
	.datad(portB31),
	.cin(gnd),
	.combout(\ShiftLeft0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~14 .lut_mask = 16'hFFF0;
defparam \ShiftLeft0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N14
cycloneive_lcell_comb \ShiftLeft0~4 (
// Equation(s):
// \ShiftLeft0~4_combout  = (\portB~41_combout ) # ((\portB~44_combout ) # ((\portB~47_combout ) # (\portB~50_combout )))

	.dataa(portB8),
	.datab(portB9),
	.datac(portB10),
	.datad(portB11),
	.cin(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~4 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N8
cycloneive_lcell_comb \ShiftLeft0~5 (
// Equation(s):
// \ShiftLeft0~5_combout  = (\portB~56_combout ) # ((\portB~62_combout ) # ((\portB~53_combout ) # (\portB~59_combout )))

	.dataa(portB13),
	.datab(portB15),
	.datac(portB12),
	.datad(portB14),
	.cin(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~5 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N20
cycloneive_lcell_comb \ShiftLeft0~3 (
// Equation(s):
// \ShiftLeft0~3_combout  = (\portB~29_combout ) # ((\portB~35_combout ) # ((\portB~38_combout ) # (\portB~32_combout )))

	.dataa(portB4),
	.datab(portB6),
	.datac(portB7),
	.datad(portB5),
	.cin(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~3 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N6
cycloneive_lcell_comb \ShiftLeft0~6 (
// Equation(s):
// \ShiftLeft0~6_combout  = (\ShiftLeft0~2_combout ) # ((\ShiftLeft0~4_combout ) # ((\ShiftLeft0~5_combout ) # (\ShiftLeft0~3_combout )))

	.dataa(\ShiftLeft0~2_combout ),
	.datab(\ShiftLeft0~4_combout ),
	.datac(\ShiftLeft0~5_combout ),
	.datad(\ShiftLeft0~3_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~6 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N16
cycloneive_lcell_comb \ShiftLeft0~7 (
// Equation(s):
// \ShiftLeft0~7_combout  = (\portB~64_combout ) # ((\portB~68_combout ) # ((\portB~66_combout ) # (\portB~70_combout )))

	.dataa(portB16),
	.datab(portB18),
	.datac(portB17),
	.datad(portB19),
	.cin(gnd),
	.combout(\ShiftLeft0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~7 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N14
cycloneive_lcell_comb \ShiftLeft0~9 (
// Equation(s):
// \ShiftLeft0~9_combout  = (\portB~87_combout ) # ((\portB~82_combout ) # (\portB~84_combout ))

	.dataa(gnd),
	.datab(portB28),
	.datac(portB26),
	.datad(portB27),
	.cin(gnd),
	.combout(\ShiftLeft0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~9 .lut_mask = 16'hFFFC;
defparam \ShiftLeft0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N0
cycloneive_lcell_comb \ShiftLeft0~11 (
// Equation(s):
// \ShiftLeft0~11_combout  = (\ShiftOp_EX~q  & (\Equal3~2_combout  & ((\portB~72_combout ) # (\portB~75_combout )))) # (!\ShiftOp_EX~q  & (((\portB~72_combout ) # (\portB~75_combout ))))

	.dataa(ShiftOp_EX),
	.datab(Equal3),
	.datac(portB20),
	.datad(portB22),
	.cin(gnd),
	.combout(\ShiftLeft0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~11 .lut_mask = 16'hDDD0;
defparam \ShiftLeft0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N6
cycloneive_lcell_comb \ShiftLeft0~12 (
// Equation(s):
// \ShiftLeft0~12_combout  = (\ShiftLeft0~8_combout ) # ((\ShiftLeft0~7_combout ) # ((\ShiftLeft0~9_combout ) # (\ShiftLeft0~11_combout )))

	.dataa(\ShiftLeft0~8_combout ),
	.datab(\ShiftLeft0~7_combout ),
	.datac(\ShiftLeft0~9_combout ),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~12 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N2
cycloneive_lcell_comb \Selector30~1 (
// Equation(s):
// \Selector30~1_combout  = (\Selector0~1_combout  & (!\portB~107_combout  & (!\ShiftLeft0~6_combout  & !\ShiftLeft0~12_combout )))

	.dataa(\Selector0~1_combout ),
	.datab(portB33),
	.datac(\ShiftLeft0~6_combout ),
	.datad(\ShiftLeft0~12_combout ),
	.cin(gnd),
	.combout(\Selector30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~1 .lut_mask = 16'h0002;
defparam \Selector30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N4
cycloneive_lcell_comb \Selector30~2 (
// Equation(s):
// \Selector30~2_combout  = (\ShiftLeft0~13_combout  & (!\portB~103_combout  & (!\ShiftLeft0~14_combout  & \Selector30~1_combout )))

	.dataa(\ShiftLeft0~13_combout ),
	.datab(portB32),
	.datac(\ShiftLeft0~14_combout ),
	.datad(\Selector30~1_combout ),
	.cin(gnd),
	.combout(\Selector30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~2 .lut_mask = 16'h0200;
defparam \Selector30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N2
cycloneive_lcell_comb \Selector0~2 (
// Equation(s):
// \Selector0~2_combout  = (ALUOp_EX[0] & (ALUOp_EX[2] & (!ALUOp_EX[3] & !ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~2 .lut_mask = 16'h0008;
defparam \Selector0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N26
cycloneive_lcell_comb \Selector30~5 (
// Equation(s):
// \Selector30~5_combout  = (Selector0 & (!\portA~12_combout  & !\portB~97_combout ))

	.dataa(Selector0),
	.datab(gnd),
	.datac(portA1),
	.datad(portB30),
	.cin(gnd),
	.combout(\Selector30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~5 .lut_mask = 16'h000A;
defparam \Selector30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N22
cycloneive_lcell_comb \Selector0~7 (
// Equation(s):
// \Selector0~7_combout  = (!ALUOp_EX[0] & (!ALUOp_EX[2] & (!ALUOp_EX[3] & ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~7 .lut_mask = 16'h0100;
defparam \Selector0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N0
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = (\portB~92_combout  & (\portA~69_combout  $ (VCC))) # (!\portB~92_combout  & (\portA~69_combout  & VCC))
// \Add0~1  = CARRY((\portB~92_combout  & \portA~69_combout ))

	.dataa(portB29),
	.datab(portA32),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h6688;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N2
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = (\portB~97_combout  & ((\portA~12_combout  & (\Add0~1  & VCC)) # (!\portA~12_combout  & (!\Add0~1 )))) # (!\portB~97_combout  & ((\portA~12_combout  & (!\Add0~1 )) # (!\portA~12_combout  & ((\Add0~1 ) # (GND)))))
// \Add0~3  = CARRY((\portB~97_combout  & (!\portA~12_combout  & !\Add0~1 )) # (!\portB~97_combout  & ((!\Add0~1 ) # (!\portA~12_combout ))))

	.dataa(portB30),
	.datab(portA1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h9617;
defparam \Add0~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N0
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (\portB~92_combout  & (\portA~69_combout  $ (VCC))) # (!\portB~92_combout  & ((\portA~69_combout ) # (GND)))
// \Add1~1  = CARRY((\portA~69_combout ) # (!\portB~92_combout ))

	.dataa(portB29),
	.datab(portA32),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h66DD;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N2
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (\portA~12_combout  & ((\portB~97_combout  & (!\Add1~1 )) # (!\portB~97_combout  & (\Add1~1  & VCC)))) # (!\portA~12_combout  & ((\portB~97_combout  & ((\Add1~1 ) # (GND))) # (!\portB~97_combout  & (!\Add1~1 ))))
// \Add1~3  = CARRY((\portA~12_combout  & (\portB~97_combout  & !\Add1~1 )) # (!\portA~12_combout  & ((\portB~97_combout ) # (!\Add1~1 ))))

	.dataa(portA1),
	.datab(portB30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h694D;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N28
cycloneive_lcell_comb \Selector30~6 (
// Equation(s):
// \Selector30~6_combout  = (\Selector0~6_combout  & ((\Add1~2_combout ) # ((\Selector0~7_combout  & \Add0~2_combout )))) # (!\Selector0~6_combout  & (\Selector0~7_combout  & (\Add0~2_combout )))

	.dataa(\Selector0~6_combout ),
	.datab(\Selector0~7_combout ),
	.datac(\Add0~2_combout ),
	.datad(\Add1~2_combout ),
	.cin(gnd),
	.combout(\Selector30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~6 .lut_mask = 16'hEAC0;
defparam \Selector30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N28
cycloneive_lcell_comb \Selector30~7 (
// Equation(s):
// \Selector30~7_combout  = (\Selector30~5_combout ) # ((\Selector30~6_combout ) # ((\Selector0~2_combout  & \portB~97_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(portB30),
	.datac(\Selector30~5_combout ),
	.datad(\Selector30~6_combout ),
	.cin(gnd),
	.combout(\Selector30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~7 .lut_mask = 16'hFFF8;
defparam \Selector30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N24
cycloneive_lcell_comb \Selector0~0 (
// Equation(s):
// \Selector0~0_combout  = (ALUOp_EX[0] & (!ALUOp_EX[2] & (!ALUOp_EX[3] & !ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~0 .lut_mask = 16'h0002;
defparam \Selector0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N26
cycloneive_lcell_comb \ShiftLeft0~8 (
// Equation(s):
// \ShiftLeft0~8_combout  = (\portB~80_combout  & (((\Equal3~2_combout )) # (!\ShiftOp_EX~q ))) # (!\portB~80_combout  & (\portB~78_combout  & ((\Equal3~2_combout ) # (!\ShiftOp_EX~q ))))

	.dataa(portB25),
	.datab(ShiftOp_EX),
	.datac(Equal3),
	.datad(portB24),
	.cin(gnd),
	.combout(\ShiftLeft0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~8 .lut_mask = 16'hF3A2;
defparam \ShiftLeft0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N24
cycloneive_lcell_comb \ShiftLeft0~10 (
// Equation(s):
// \ShiftLeft0~10_combout  = (\portB~76_combout ) # ((\portB~73_combout ) # ((\ShiftLeft0~8_combout ) # (\ShiftLeft0~9_combout )))

	.dataa(portB23),
	.datab(portB21),
	.datac(\ShiftLeft0~8_combout ),
	.datad(\ShiftLeft0~9_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~10 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N28
cycloneive_lcell_comb \Selector31~0 (
// Equation(s):
// \Selector31~0_combout  = (!\ShiftLeft0~7_combout  & (\Selector0~0_combout  & (!\ShiftLeft0~6_combout  & !\ShiftLeft0~10_combout )))

	.dataa(\ShiftLeft0~7_combout ),
	.datab(\Selector0~0_combout ),
	.datac(\ShiftLeft0~6_combout ),
	.datad(\ShiftLeft0~10_combout ),
	.cin(gnd),
	.combout(\Selector31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~0 .lut_mask = 16'h0004;
defparam \Selector31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N2
cycloneive_lcell_comb \ShiftRight0~13 (
// Equation(s):
// \ShiftRight0~13_combout  = (\portB~92_combout  & (\portA~36_combout )) # (!\portB~92_combout  & ((\portA~37_combout )))

	.dataa(gnd),
	.datab(portA15),
	.datac(portA16),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~13 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N16
cycloneive_lcell_comb \ShiftRight0~12 (
// Equation(s):
// \ShiftRight0~12_combout  = (\portB~92_combout  & ((\portA~33_combout ))) # (!\portB~92_combout  & (\portA~35_combout ))

	.dataa(portA14),
	.datab(gnd),
	.datac(portA13),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~12 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N28
cycloneive_lcell_comb \ShiftRight0~14 (
// Equation(s):
// \ShiftRight0~14_combout  = (\portB~97_combout  & ((\ShiftRight0~12_combout ))) # (!\portB~97_combout  & (\ShiftRight0~13_combout ))

	.dataa(portB30),
	.datab(\ShiftRight0~13_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~12_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~14 .lut_mask = 16'hEE44;
defparam \ShiftRight0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N18
cycloneive_lcell_comb \ShiftRight0~15 (
// Equation(s):
// \ShiftRight0~15_combout  = (\portB~100_combout  & (\ShiftRight0~11_combout )) # (!\portB~100_combout  & ((\ShiftRight0~14_combout )))

	.dataa(\ShiftRight0~11_combout ),
	.datab(portB31),
	.datac(gnd),
	.datad(\ShiftRight0~14_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~15 .lut_mask = 16'hBB88;
defparam \ShiftRight0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N24
cycloneive_lcell_comb \ShiftRight0~6 (
// Equation(s):
// \ShiftRight0~6_combout  = (\portB~92_combout  & (\portA~21_combout )) # (!\portB~92_combout  & ((\portA~23_combout )))

	.dataa(gnd),
	.datab(portA7),
	.datac(portA8),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~6 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N14
cycloneive_lcell_comb \ShiftRight0~5 (
// Equation(s):
// \ShiftRight0~5_combout  = (\portB~92_combout  & (\portA~17_combout )) # (!\portB~92_combout  & ((\portA~19_combout )))

	.dataa(gnd),
	.datab(portA5),
	.datac(portA6),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~5 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N14
cycloneive_lcell_comb \ShiftRight0~7 (
// Equation(s):
// \ShiftRight0~7_combout  = (\portB~97_combout  & ((\ShiftRight0~5_combout ))) # (!\portB~97_combout  & (\ShiftRight0~6_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~6_combout ),
	.datac(portB30),
	.datad(\ShiftRight0~5_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~7 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N28
cycloneive_lcell_comb \ShiftRight0~3 (
// Equation(s):
// \ShiftRight0~3_combout  = (\portB~92_combout  & ((\portA~14_combout ))) # (!\portB~92_combout  & (\portA~16_combout ))

	.dataa(portA4),
	.datab(portA2),
	.datac(gnd),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~3_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~3 .lut_mask = 16'hCCAA;
defparam \ShiftRight0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N22
cycloneive_lcell_comb \ShiftRight0~2 (
// Equation(s):
// \ShiftRight0~2_combout  = (!\portB~97_combout  & ((\portB~92_combout  & (\portA~9_combout )) # (!\portB~92_combout  & ((\portA~12_combout )))))

	.dataa(portB29),
	.datab(portA),
	.datac(portA1),
	.datad(portB30),
	.cin(gnd),
	.combout(\ShiftRight0~2_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~2 .lut_mask = 16'h00D8;
defparam \ShiftRight0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N12
cycloneive_lcell_comb \ShiftRight0~4 (
// Equation(s):
// \ShiftRight0~4_combout  = (!\portB~100_combout  & ((\ShiftRight0~2_combout ) # ((\ShiftRight0~3_combout  & \portB~97_combout ))))

	.dataa(portB31),
	.datab(\ShiftRight0~3_combout ),
	.datac(\ShiftRight0~2_combout ),
	.datad(portB30),
	.cin(gnd),
	.combout(\ShiftRight0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~4 .lut_mask = 16'h5450;
defparam \ShiftRight0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N12
cycloneive_lcell_comb \ShiftRight0~8 (
// Equation(s):
// \ShiftRight0~8_combout  = (!\portB~103_combout  & ((\ShiftRight0~4_combout ) # ((\portB~100_combout  & \ShiftRight0~7_combout ))))

	.dataa(portB31),
	.datab(portB32),
	.datac(\ShiftRight0~7_combout ),
	.datad(\ShiftRight0~4_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~8 .lut_mask = 16'h3320;
defparam \ShiftRight0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N14
cycloneive_lcell_comb \ShiftRight0~16 (
// Equation(s):
// \ShiftRight0~16_combout  = (!\portB~107_combout  & ((\ShiftRight0~8_combout ) # ((\portB~103_combout  & \ShiftRight0~15_combout ))))

	.dataa(portB33),
	.datab(portB32),
	.datac(\ShiftRight0~15_combout ),
	.datad(\ShiftRight0~8_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~16 .lut_mask = 16'h5540;
defparam \ShiftRight0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N28
cycloneive_lcell_comb \ShiftRight0~20 (
// Equation(s):
// \ShiftRight0~20_combout  = (\portB~92_combout  & (\portA~49_combout )) # (!\portB~92_combout  & ((\portA~51_combout )))

	.dataa(portA22),
	.datab(gnd),
	.datac(portA23),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~20 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N24
cycloneive_lcell_comb \ShiftRight0~19 (
// Equation(s):
// \ShiftRight0~19_combout  = (\portB~92_combout  & ((\portA~45_combout ))) # (!\portB~92_combout  & (\portA~47_combout ))

	.dataa(portA21),
	.datab(gnd),
	.datac(portB29),
	.datad(portA20),
	.cin(gnd),
	.combout(\ShiftRight0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~19 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N4
cycloneive_lcell_comb \ShiftRight0~21 (
// Equation(s):
// \ShiftRight0~21_combout  = (\portB~97_combout  & ((\ShiftRight0~19_combout ))) # (!\portB~97_combout  & (\ShiftRight0~20_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftRight0~20_combout ),
	.datad(\ShiftRight0~19_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~21 .lut_mask = 16'hFA50;
defparam \ShiftRight0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N20
cycloneive_lcell_comb \ShiftRight0~17 (
// Equation(s):
// \ShiftRight0~17_combout  = (!\portB~92_combout  & ((\portB~97_combout  & ((\portA~39_combout ))) # (!\portB~97_combout  & (\portA~41_combout ))))

	.dataa(portA18),
	.datab(portB30),
	.datac(portA17),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~17 .lut_mask = 16'h00E2;
defparam \ShiftRight0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N2
cycloneive_lcell_comb \ShiftRight0~18 (
// Equation(s):
// \ShiftRight0~18_combout  = (\ShiftRight0~17_combout ) # ((\portB~92_combout  & (\portA~43_combout  & !\portB~97_combout )))

	.dataa(portB29),
	.datab(portA19),
	.datac(portB30),
	.datad(\ShiftRight0~17_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~18 .lut_mask = 16'hFF08;
defparam \ShiftRight0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N6
cycloneive_lcell_comb \ShiftRight0~22 (
// Equation(s):
// \ShiftRight0~22_combout  = (\portB~100_combout  & ((\ShiftRight0~18_combout ))) # (!\portB~100_combout  & (\ShiftRight0~21_combout ))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftRight0~21_combout ),
	.datad(\ShiftRight0~18_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~22 .lut_mask = 16'hFC30;
defparam \ShiftRight0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N12
cycloneive_lcell_comb \ShiftRight0~26 (
// Equation(s):
// \ShiftRight0~26_combout  = (\portB~92_combout  & (\portA~61_combout )) # (!\portB~92_combout  & ((\portA~63_combout )))

	.dataa(portA28),
	.datab(gnd),
	.datac(portA29),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~26 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N6
cycloneive_lcell_comb \ShiftRight0~27 (
// Equation(s):
// \ShiftRight0~27_combout  = (\portB~92_combout  & (\portA~65_combout )) # (!\portB~92_combout  & ((\portA~67_combout )))

	.dataa(portA30),
	.datab(gnd),
	.datac(portA31),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~27 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N26
cycloneive_lcell_comb \ShiftRight0~28 (
// Equation(s):
// \ShiftRight0~28_combout  = (\portB~97_combout  & (\ShiftRight0~26_combout )) # (!\portB~97_combout  & ((\ShiftRight0~27_combout )))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftRight0~26_combout ),
	.datad(\ShiftRight0~27_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~28 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N30
cycloneive_lcell_comb \ShiftRight0~24 (
// Equation(s):
// \ShiftRight0~24_combout  = (\portB~92_combout  & ((\portA~57_combout ))) # (!\portB~92_combout  & (\portA~59_combout ))

	.dataa(portA27),
	.datab(gnd),
	.datac(portA26),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~24 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N14
cycloneive_lcell_comb \ShiftRight0~23 (
// Equation(s):
// \ShiftRight0~23_combout  = (\portB~92_combout  & ((\portA~53_combout ))) # (!\portB~92_combout  & (\portA~55_combout ))

	.dataa(gnd),
	.datab(portA25),
	.datac(portA24),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~23 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N20
cycloneive_lcell_comb \ShiftRight0~25 (
// Equation(s):
// \ShiftRight0~25_combout  = (\portB~97_combout  & ((\ShiftRight0~23_combout ))) # (!\portB~97_combout  & (\ShiftRight0~24_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftRight0~24_combout ),
	.datad(\ShiftRight0~23_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~25 .lut_mask = 16'hFA50;
defparam \ShiftRight0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N28
cycloneive_lcell_comb \Selector22~0 (
// Equation(s):
// \Selector22~0_combout  = (\portB~100_combout  & ((\ShiftRight0~25_combout ))) # (!\portB~100_combout  & (\ShiftRight0~28_combout ))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftRight0~28_combout ),
	.datad(\ShiftRight0~25_combout ),
	.cin(gnd),
	.combout(\Selector22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~0 .lut_mask = 16'hFC30;
defparam \Selector22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N12
cycloneive_lcell_comb \ShiftRight0~29 (
// Equation(s):
// \ShiftRight0~29_combout  = (\portB~103_combout  & (\ShiftRight0~22_combout )) # (!\portB~103_combout  & ((\Selector22~0_combout )))

	.dataa(portB32),
	.datab(gnd),
	.datac(\ShiftRight0~22_combout ),
	.datad(\Selector22~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~29 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N28
cycloneive_lcell_comb \Selector30~0 (
// Equation(s):
// \Selector30~0_combout  = (\Selector31~0_combout  & ((\ShiftRight0~16_combout ) # ((\portB~107_combout  & \ShiftRight0~29_combout ))))

	.dataa(portB33),
	.datab(\Selector31~0_combout ),
	.datac(\ShiftRight0~16_combout ),
	.datad(\ShiftRight0~29_combout ),
	.cin(gnd),
	.combout(\Selector30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~0 .lut_mask = 16'hC8C0;
defparam \Selector30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N16
cycloneive_lcell_comb \Selector0~6 (
// Equation(s):
// \Selector0~6_combout  = (ALUOp_EX[0] & (!ALUOp_EX[2] & (!ALUOp_EX[3] & ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~6 .lut_mask = 16'h0200;
defparam \Selector0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N18
cycloneive_lcell_comb \Selector31~2 (
// Equation(s):
// \Selector31~2_combout  = (\Selector0~2_combout  & ((\portB~92_combout ) # ((\Selector0~6_combout  & \Add1~0_combout )))) # (!\Selector0~2_combout  & (\Selector0~6_combout  & (\Add1~0_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(\Selector0~6_combout ),
	.datac(\Add1~0_combout ),
	.datad(portB29),
	.cin(gnd),
	.combout(\Selector31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~2 .lut_mask = 16'hEAC0;
defparam \Selector31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N4
cycloneive_lcell_comb \Selector31~3 (
// Equation(s):
// \Selector31~3_combout  = (\Selector31~2_combout ) # ((\Add0~0_combout  & ((\Selector0~4_combout ) # (\Selector0~7_combout ))))

	.dataa(\Selector0~4_combout ),
	.datab(\Selector0~7_combout ),
	.datac(\Add0~0_combout ),
	.datad(\Selector31~2_combout ),
	.cin(gnd),
	.combout(\Selector31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~3 .lut_mask = 16'hFFE0;
defparam \Selector31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N0
cycloneive_lcell_comb \LessThan1~1 (
// Equation(s):
// \LessThan1~1_cout  = CARRY((\portB~92_combout  & !\portA~69_combout ))

	.dataa(portB29),
	.datab(portA32),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan1~1_cout ));
// synopsys translate_off
defparam \LessThan1~1 .lut_mask = 16'h0022;
defparam \LessThan1~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N2
cycloneive_lcell_comb \LessThan1~3 (
// Equation(s):
// \LessThan1~3_cout  = CARRY((\portA~12_combout  & ((!\LessThan1~1_cout ) # (!\portB~97_combout ))) # (!\portA~12_combout  & (!\portB~97_combout  & !\LessThan1~1_cout )))

	.dataa(portA1),
	.datab(portB30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~1_cout ),
	.combout(),
	.cout(\LessThan1~3_cout ));
// synopsys translate_off
defparam \LessThan1~3 .lut_mask = 16'h002B;
defparam \LessThan1~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N4
cycloneive_lcell_comb \LessThan1~5 (
// Equation(s):
// \LessThan1~5_cout  = CARRY((\portA~9_combout  & (\portB~100_combout  & !\LessThan1~3_cout )) # (!\portA~9_combout  & ((\portB~100_combout ) # (!\LessThan1~3_cout ))))

	.dataa(portA),
	.datab(portB31),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~3_cout ),
	.combout(),
	.cout(\LessThan1~5_cout ));
// synopsys translate_off
defparam \LessThan1~5 .lut_mask = 16'h004D;
defparam \LessThan1~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N6
cycloneive_lcell_comb \LessThan1~7 (
// Equation(s):
// \LessThan1~7_cout  = CARRY((\portA~16_combout  & ((!\LessThan1~5_cout ) # (!\portB~103_combout ))) # (!\portA~16_combout  & (!\portB~103_combout  & !\LessThan1~5_cout )))

	.dataa(portA4),
	.datab(portB32),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~5_cout ),
	.combout(),
	.cout(\LessThan1~7_cout ));
// synopsys translate_off
defparam \LessThan1~7 .lut_mask = 16'h002B;
defparam \LessThan1~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N8
cycloneive_lcell_comb \LessThan1~9 (
// Equation(s):
// \LessThan1~9_cout  = CARRY((\portA~14_combout  & (\portB~107_combout  & !\LessThan1~7_cout )) # (!\portA~14_combout  & ((\portB~107_combout ) # (!\LessThan1~7_cout ))))

	.dataa(portA2),
	.datab(portB33),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~7_cout ),
	.combout(),
	.cout(\LessThan1~9_cout ));
// synopsys translate_off
defparam \LessThan1~9 .lut_mask = 16'h004D;
defparam \LessThan1~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N10
cycloneive_lcell_comb \LessThan1~11 (
// Equation(s):
// \LessThan1~11_cout  = CARRY((\portB~87_combout  & (\portA~23_combout  & !\LessThan1~9_cout )) # (!\portB~87_combout  & ((\portA~23_combout ) # (!\LessThan1~9_cout ))))

	.dataa(portB28),
	.datab(portA8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~9_cout ),
	.combout(),
	.cout(\LessThan1~11_cout ));
// synopsys translate_off
defparam \LessThan1~11 .lut_mask = 16'h004D;
defparam \LessThan1~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N12
cycloneive_lcell_comb \LessThan1~13 (
// Equation(s):
// \LessThan1~13_cout  = CARRY((\portA~21_combout  & (\portB~84_combout  & !\LessThan1~11_cout )) # (!\portA~21_combout  & ((\portB~84_combout ) # (!\LessThan1~11_cout ))))

	.dataa(portA7),
	.datab(portB27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~11_cout ),
	.combout(),
	.cout(\LessThan1~13_cout ));
// synopsys translate_off
defparam \LessThan1~13 .lut_mask = 16'h004D;
defparam \LessThan1~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N14
cycloneive_lcell_comb \LessThan1~15 (
// Equation(s):
// \LessThan1~15_cout  = CARRY((\portB~82_combout  & (\portA~19_combout  & !\LessThan1~13_cout )) # (!\portB~82_combout  & ((\portA~19_combout ) # (!\LessThan1~13_cout ))))

	.dataa(portB26),
	.datab(portA6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~13_cout ),
	.combout(),
	.cout(\LessThan1~15_cout ));
// synopsys translate_off
defparam \LessThan1~15 .lut_mask = 16'h004D;
defparam \LessThan1~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N16
cycloneive_lcell_comb \LessThan1~17 (
// Equation(s):
// \LessThan1~17_cout  = CARRY((\portB~76_combout  & ((!\LessThan1~15_cout ) # (!\portA~17_combout ))) # (!\portB~76_combout  & (!\portA~17_combout  & !\LessThan1~15_cout )))

	.dataa(portB23),
	.datab(portA5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~15_cout ),
	.combout(),
	.cout(\LessThan1~17_cout ));
// synopsys translate_off
defparam \LessThan1~17 .lut_mask = 16'h002B;
defparam \LessThan1~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N18
cycloneive_lcell_comb \LessThan1~19 (
// Equation(s):
// \LessThan1~19_cout  = CARRY((\portA~37_combout  & ((!\LessThan1~17_cout ) # (!\portB~73_combout ))) # (!\portA~37_combout  & (!\portB~73_combout  & !\LessThan1~17_cout )))

	.dataa(portA16),
	.datab(portB21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~17_cout ),
	.combout(),
	.cout(\LessThan1~19_cout ));
// synopsys translate_off
defparam \LessThan1~19 .lut_mask = 16'h002B;
defparam \LessThan1~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N20
cycloneive_lcell_comb \LessThan1~21 (
// Equation(s):
// \LessThan1~21_cout  = CARRY((\portB~109_combout  & ((!\LessThan1~19_cout ) # (!\portA~36_combout ))) # (!\portB~109_combout  & (!\portA~36_combout  & !\LessThan1~19_cout )))

	.dataa(portB35),
	.datab(portA15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~19_cout ),
	.combout(),
	.cout(\LessThan1~21_cout ));
// synopsys translate_off
defparam \LessThan1~21 .lut_mask = 16'h002B;
defparam \LessThan1~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N22
cycloneive_lcell_comb \LessThan1~23 (
// Equation(s):
// \LessThan1~23_cout  = CARRY((\portB~108_combout  & (\portA~35_combout  & !\LessThan1~21_cout )) # (!\portB~108_combout  & ((\portA~35_combout ) # (!\LessThan1~21_cout ))))

	.dataa(portB34),
	.datab(portA14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~21_cout ),
	.combout(),
	.cout(\LessThan1~23_cout ));
// synopsys translate_off
defparam \LessThan1~23 .lut_mask = 16'h004D;
defparam \LessThan1~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N24
cycloneive_lcell_comb \LessThan1~25 (
// Equation(s):
// \LessThan1~25_cout  = CARRY((\portB~70_combout  & ((!\LessThan1~23_cout ) # (!\portA~33_combout ))) # (!\portB~70_combout  & (!\portA~33_combout  & !\LessThan1~23_cout )))

	.dataa(portB19),
	.datab(portA13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~23_cout ),
	.combout(),
	.cout(\LessThan1~25_cout ));
// synopsys translate_off
defparam \LessThan1~25 .lut_mask = 16'h002B;
defparam \LessThan1~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N26
cycloneive_lcell_comb \LessThan1~27 (
// Equation(s):
// \LessThan1~27_cout  = CARRY((\portB~68_combout  & (\portA~31_combout  & !\LessThan1~25_cout )) # (!\portB~68_combout  & ((\portA~31_combout ) # (!\LessThan1~25_cout ))))

	.dataa(portB18),
	.datab(portA12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~25_cout ),
	.combout(),
	.cout(\LessThan1~27_cout ));
// synopsys translate_off
defparam \LessThan1~27 .lut_mask = 16'h004D;
defparam \LessThan1~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N28
cycloneive_lcell_comb \LessThan1~29 (
// Equation(s):
// \LessThan1~29_cout  = CARRY((\portA~29_combout  & (\portB~66_combout  & !\LessThan1~27_cout )) # (!\portA~29_combout  & ((\portB~66_combout ) # (!\LessThan1~27_cout ))))

	.dataa(portA11),
	.datab(portB17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~27_cout ),
	.combout(),
	.cout(\LessThan1~29_cout ));
// synopsys translate_off
defparam \LessThan1~29 .lut_mask = 16'h004D;
defparam \LessThan1~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N30
cycloneive_lcell_comb \LessThan1~31 (
// Equation(s):
// \LessThan1~31_cout  = CARRY((\portB~64_combout  & (\portA~27_combout  & !\LessThan1~29_cout )) # (!\portB~64_combout  & ((\portA~27_combout ) # (!\LessThan1~29_cout ))))

	.dataa(portB16),
	.datab(portA10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~29_cout ),
	.combout(),
	.cout(\LessThan1~31_cout ));
// synopsys translate_off
defparam \LessThan1~31 .lut_mask = 16'h004D;
defparam \LessThan1~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N0
cycloneive_lcell_comb \LessThan1~33 (
// Equation(s):
// \LessThan1~33_cout  = CARRY((\portB~62_combout  & ((!\LessThan1~31_cout ) # (!\portA~25_combout ))) # (!\portB~62_combout  & (!\portA~25_combout  & !\LessThan1~31_cout )))

	.dataa(portB15),
	.datab(portA9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~31_cout ),
	.combout(),
	.cout(\LessThan1~33_cout ));
// synopsys translate_off
defparam \LessThan1~33 .lut_mask = 16'h002B;
defparam \LessThan1~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N2
cycloneive_lcell_comb \LessThan1~35 (
// Equation(s):
// \LessThan1~35_cout  = CARRY((\portB~59_combout  & (\portA~67_combout  & !\LessThan1~33_cout )) # (!\portB~59_combout  & ((\portA~67_combout ) # (!\LessThan1~33_cout ))))

	.dataa(portB14),
	.datab(portA31),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~33_cout ),
	.combout(),
	.cout(\LessThan1~35_cout ));
// synopsys translate_off
defparam \LessThan1~35 .lut_mask = 16'h004D;
defparam \LessThan1~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N4
cycloneive_lcell_comb \LessThan1~37 (
// Equation(s):
// \LessThan1~37_cout  = CARRY((\portB~56_combout  & ((!\LessThan1~35_cout ) # (!\portA~65_combout ))) # (!\portB~56_combout  & (!\portA~65_combout  & !\LessThan1~35_cout )))

	.dataa(portB13),
	.datab(portA30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~35_cout ),
	.combout(),
	.cout(\LessThan1~37_cout ));
// synopsys translate_off
defparam \LessThan1~37 .lut_mask = 16'h002B;
defparam \LessThan1~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N6
cycloneive_lcell_comb \LessThan1~39 (
// Equation(s):
// \LessThan1~39_cout  = CARRY((\portA~63_combout  & ((!\LessThan1~37_cout ) # (!\portB~53_combout ))) # (!\portA~63_combout  & (!\portB~53_combout  & !\LessThan1~37_cout )))

	.dataa(portA29),
	.datab(portB12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~37_cout ),
	.combout(),
	.cout(\LessThan1~39_cout ));
// synopsys translate_off
defparam \LessThan1~39 .lut_mask = 16'h002B;
defparam \LessThan1~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N8
cycloneive_lcell_comb \LessThan1~41 (
// Equation(s):
// \LessThan1~41_cout  = CARRY((\portA~61_combout  & (\portB~50_combout  & !\LessThan1~39_cout )) # (!\portA~61_combout  & ((\portB~50_combout ) # (!\LessThan1~39_cout ))))

	.dataa(portA28),
	.datab(portB11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~39_cout ),
	.combout(),
	.cout(\LessThan1~41_cout ));
// synopsys translate_off
defparam \LessThan1~41 .lut_mask = 16'h004D;
defparam \LessThan1~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N10
cycloneive_lcell_comb \LessThan1~43 (
// Equation(s):
// \LessThan1~43_cout  = CARRY((\portA~59_combout  & ((!\LessThan1~41_cout ) # (!\portB~47_combout ))) # (!\portA~59_combout  & (!\portB~47_combout  & !\LessThan1~41_cout )))

	.dataa(portA27),
	.datab(portB10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~41_cout ),
	.combout(),
	.cout(\LessThan1~43_cout ));
// synopsys translate_off
defparam \LessThan1~43 .lut_mask = 16'h002B;
defparam \LessThan1~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N12
cycloneive_lcell_comb \LessThan1~45 (
// Equation(s):
// \LessThan1~45_cout  = CARRY((\portB~44_combout  & ((!\LessThan1~43_cout ) # (!\portA~57_combout ))) # (!\portB~44_combout  & (!\portA~57_combout  & !\LessThan1~43_cout )))

	.dataa(portB9),
	.datab(portA26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~43_cout ),
	.combout(),
	.cout(\LessThan1~45_cout ));
// synopsys translate_off
defparam \LessThan1~45 .lut_mask = 16'h002B;
defparam \LessThan1~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N14
cycloneive_lcell_comb \LessThan1~47 (
// Equation(s):
// \LessThan1~47_cout  = CARRY((\portB~41_combout  & (\portA~55_combout  & !\LessThan1~45_cout )) # (!\portB~41_combout  & ((\portA~55_combout ) # (!\LessThan1~45_cout ))))

	.dataa(portB8),
	.datab(portA25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~45_cout ),
	.combout(),
	.cout(\LessThan1~47_cout ));
// synopsys translate_off
defparam \LessThan1~47 .lut_mask = 16'h004D;
defparam \LessThan1~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N16
cycloneive_lcell_comb \LessThan1~49 (
// Equation(s):
// \LessThan1~49_cout  = CARRY((\portB~38_combout  & ((!\LessThan1~47_cout ) # (!\portA~53_combout ))) # (!\portB~38_combout  & (!\portA~53_combout  & !\LessThan1~47_cout )))

	.dataa(portB7),
	.datab(portA24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~47_cout ),
	.combout(),
	.cout(\LessThan1~49_cout ));
// synopsys translate_off
defparam \LessThan1~49 .lut_mask = 16'h002B;
defparam \LessThan1~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N18
cycloneive_lcell_comb \LessThan1~51 (
// Equation(s):
// \LessThan1~51_cout  = CARRY((\portB~35_combout  & (\portA~51_combout  & !\LessThan1~49_cout )) # (!\portB~35_combout  & ((\portA~51_combout ) # (!\LessThan1~49_cout ))))

	.dataa(portB6),
	.datab(portA23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~49_cout ),
	.combout(),
	.cout(\LessThan1~51_cout ));
// synopsys translate_off
defparam \LessThan1~51 .lut_mask = 16'h004D;
defparam \LessThan1~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N20
cycloneive_lcell_comb \LessThan1~53 (
// Equation(s):
// \LessThan1~53_cout  = CARRY((\portB~32_combout  & ((!\LessThan1~51_cout ) # (!\portA~49_combout ))) # (!\portB~32_combout  & (!\portA~49_combout  & !\LessThan1~51_cout )))

	.dataa(portB5),
	.datab(portA22),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~51_cout ),
	.combout(),
	.cout(\LessThan1~53_cout ));
// synopsys translate_off
defparam \LessThan1~53 .lut_mask = 16'h002B;
defparam \LessThan1~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N22
cycloneive_lcell_comb \LessThan1~55 (
// Equation(s):
// \LessThan1~55_cout  = CARRY((\portB~29_combout  & (\portA~47_combout  & !\LessThan1~53_cout )) # (!\portB~29_combout  & ((\portA~47_combout ) # (!\LessThan1~53_cout ))))

	.dataa(portB4),
	.datab(portA21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~53_cout ),
	.combout(),
	.cout(\LessThan1~55_cout ));
// synopsys translate_off
defparam \LessThan1~55 .lut_mask = 16'h004D;
defparam \LessThan1~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N24
cycloneive_lcell_comb \LessThan1~57 (
// Equation(s):
// \LessThan1~57_cout  = CARRY((\portB~26_combout  & ((!\LessThan1~55_cout ) # (!\portA~45_combout ))) # (!\portB~26_combout  & (!\portA~45_combout  & !\LessThan1~55_cout )))

	.dataa(portB3),
	.datab(portA20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~55_cout ),
	.combout(),
	.cout(\LessThan1~57_cout ));
// synopsys translate_off
defparam \LessThan1~57 .lut_mask = 16'h002B;
defparam \LessThan1~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N26
cycloneive_lcell_comb \LessThan1~59 (
// Equation(s):
// \LessThan1~59_cout  = CARRY((\portA~41_combout  & ((!\LessThan1~57_cout ) # (!\portB~23_combout ))) # (!\portA~41_combout  & (!\portB~23_combout  & !\LessThan1~57_cout )))

	.dataa(portA18),
	.datab(portB2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~57_cout ),
	.combout(),
	.cout(\LessThan1~59_cout ));
// synopsys translate_off
defparam \LessThan1~59 .lut_mask = 16'h002B;
defparam \LessThan1~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N28
cycloneive_lcell_comb \LessThan1~61 (
// Equation(s):
// \LessThan1~61_cout  = CARRY((\portA~43_combout  & (\portB~20_combout  & !\LessThan1~59_cout )) # (!\portA~43_combout  & ((\portB~20_combout ) # (!\LessThan1~59_cout ))))

	.dataa(portA19),
	.datab(portB1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~59_cout ),
	.combout(),
	.cout(\LessThan1~61_cout ));
// synopsys translate_off
defparam \LessThan1~61 .lut_mask = 16'h004D;
defparam \LessThan1~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N30
cycloneive_lcell_comb \LessThan1~62 (
// Equation(s):
// \LessThan1~62_combout  = (\portA~39_combout  & (\LessThan1~61_cout  & \portB~17_combout )) # (!\portA~39_combout  & ((\LessThan1~61_cout ) # (\portB~17_combout )))

	.dataa(gnd),
	.datab(portA17),
	.datac(gnd),
	.datad(portB),
	.cin(\LessThan1~61_cout ),
	.combout(\LessThan1~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~62 .lut_mask = 16'hF330;
defparam \LessThan1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N0
cycloneive_lcell_comb \LessThan0~1 (
// Equation(s):
// \LessThan0~1_cout  = CARRY((!\portA~69_combout  & \portB~92_combout ))

	.dataa(portA32),
	.datab(portB29),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
// synopsys translate_off
defparam \LessThan0~1 .lut_mask = 16'h0044;
defparam \LessThan0~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N2
cycloneive_lcell_comb \LessThan0~3 (
// Equation(s):
// \LessThan0~3_cout  = CARRY((\portA~12_combout  & ((!\LessThan0~1_cout ) # (!\portB~97_combout ))) # (!\portA~12_combout  & (!\portB~97_combout  & !\LessThan0~1_cout )))

	.dataa(portA1),
	.datab(portB30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
// synopsys translate_off
defparam \LessThan0~3 .lut_mask = 16'h002B;
defparam \LessThan0~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N4
cycloneive_lcell_comb \LessThan0~5 (
// Equation(s):
// \LessThan0~5_cout  = CARRY((\portB~100_combout  & ((!\LessThan0~3_cout ) # (!\portA~9_combout ))) # (!\portB~100_combout  & (!\portA~9_combout  & !\LessThan0~3_cout )))

	.dataa(portB31),
	.datab(portA),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
// synopsys translate_off
defparam \LessThan0~5 .lut_mask = 16'h002B;
defparam \LessThan0~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N6
cycloneive_lcell_comb \LessThan0~7 (
// Equation(s):
// \LessThan0~7_cout  = CARRY((\portA~16_combout  & ((!\LessThan0~5_cout ) # (!\portB~103_combout ))) # (!\portA~16_combout  & (!\portB~103_combout  & !\LessThan0~5_cout )))

	.dataa(portA4),
	.datab(portB32),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
// synopsys translate_off
defparam \LessThan0~7 .lut_mask = 16'h002B;
defparam \LessThan0~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N8
cycloneive_lcell_comb \LessThan0~9 (
// Equation(s):
// \LessThan0~9_cout  = CARRY((\portA~14_combout  & (\portB~107_combout  & !\LessThan0~7_cout )) # (!\portA~14_combout  & ((\portB~107_combout ) # (!\LessThan0~7_cout ))))

	.dataa(portA2),
	.datab(portB33),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
// synopsys translate_off
defparam \LessThan0~9 .lut_mask = 16'h004D;
defparam \LessThan0~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N10
cycloneive_lcell_comb \LessThan0~11 (
// Equation(s):
// \LessThan0~11_cout  = CARRY((\portA~23_combout  & ((!\LessThan0~9_cout ) # (!\portB~87_combout ))) # (!\portA~23_combout  & (!\portB~87_combout  & !\LessThan0~9_cout )))

	.dataa(portA8),
	.datab(portB28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
// synopsys translate_off
defparam \LessThan0~11 .lut_mask = 16'h002B;
defparam \LessThan0~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N12
cycloneive_lcell_comb \LessThan0~13 (
// Equation(s):
// \LessThan0~13_cout  = CARRY((\portB~84_combout  & ((!\LessThan0~11_cout ) # (!\portA~21_combout ))) # (!\portB~84_combout  & (!\portA~21_combout  & !\LessThan0~11_cout )))

	.dataa(portB27),
	.datab(portA7),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
// synopsys translate_off
defparam \LessThan0~13 .lut_mask = 16'h002B;
defparam \LessThan0~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N14
cycloneive_lcell_comb \LessThan0~15 (
// Equation(s):
// \LessThan0~15_cout  = CARRY((\portB~82_combout  & (\portA~19_combout  & !\LessThan0~13_cout )) # (!\portB~82_combout  & ((\portA~19_combout ) # (!\LessThan0~13_cout ))))

	.dataa(portB26),
	.datab(portA6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
// synopsys translate_off
defparam \LessThan0~15 .lut_mask = 16'h004D;
defparam \LessThan0~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N16
cycloneive_lcell_comb \LessThan0~17 (
// Equation(s):
// \LessThan0~17_cout  = CARRY((\portA~17_combout  & (\portB~76_combout  & !\LessThan0~15_cout )) # (!\portA~17_combout  & ((\portB~76_combout ) # (!\LessThan0~15_cout ))))

	.dataa(portA5),
	.datab(portB23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
// synopsys translate_off
defparam \LessThan0~17 .lut_mask = 16'h004D;
defparam \LessThan0~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N18
cycloneive_lcell_comb \LessThan0~19 (
// Equation(s):
// \LessThan0~19_cout  = CARRY((\portA~37_combout  & ((!\LessThan0~17_cout ) # (!\portB~73_combout ))) # (!\portA~37_combout  & (!\portB~73_combout  & !\LessThan0~17_cout )))

	.dataa(portA16),
	.datab(portB21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
// synopsys translate_off
defparam \LessThan0~19 .lut_mask = 16'h002B;
defparam \LessThan0~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N20
cycloneive_lcell_comb \LessThan0~21 (
// Equation(s):
// \LessThan0~21_cout  = CARRY((\portB~109_combout  & ((!\LessThan0~19_cout ) # (!\portA~36_combout ))) # (!\portB~109_combout  & (!\portA~36_combout  & !\LessThan0~19_cout )))

	.dataa(portB35),
	.datab(portA15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
// synopsys translate_off
defparam \LessThan0~21 .lut_mask = 16'h002B;
defparam \LessThan0~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N22
cycloneive_lcell_comb \LessThan0~23 (
// Equation(s):
// \LessThan0~23_cout  = CARRY((\portA~35_combout  & ((!\LessThan0~21_cout ) # (!\portB~108_combout ))) # (!\portA~35_combout  & (!\portB~108_combout  & !\LessThan0~21_cout )))

	.dataa(portA14),
	.datab(portB34),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~21_cout ),
	.combout(),
	.cout(\LessThan0~23_cout ));
// synopsys translate_off
defparam \LessThan0~23 .lut_mask = 16'h002B;
defparam \LessThan0~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N24
cycloneive_lcell_comb \LessThan0~25 (
// Equation(s):
// \LessThan0~25_cout  = CARRY((\portB~70_combout  & ((!\LessThan0~23_cout ) # (!\portA~33_combout ))) # (!\portB~70_combout  & (!\portA~33_combout  & !\LessThan0~23_cout )))

	.dataa(portB19),
	.datab(portA13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~23_cout ),
	.combout(),
	.cout(\LessThan0~25_cout ));
// synopsys translate_off
defparam \LessThan0~25 .lut_mask = 16'h002B;
defparam \LessThan0~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N26
cycloneive_lcell_comb \LessThan0~27 (
// Equation(s):
// \LessThan0~27_cout  = CARRY((\portA~31_combout  & ((!\LessThan0~25_cout ) # (!\portB~68_combout ))) # (!\portA~31_combout  & (!\portB~68_combout  & !\LessThan0~25_cout )))

	.dataa(portA12),
	.datab(portB18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~25_cout ),
	.combout(),
	.cout(\LessThan0~27_cout ));
// synopsys translate_off
defparam \LessThan0~27 .lut_mask = 16'h002B;
defparam \LessThan0~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N28
cycloneive_lcell_comb \LessThan0~29 (
// Equation(s):
// \LessThan0~29_cout  = CARRY((\portB~66_combout  & ((!\LessThan0~27_cout ) # (!\portA~29_combout ))) # (!\portB~66_combout  & (!\portA~29_combout  & !\LessThan0~27_cout )))

	.dataa(portB17),
	.datab(portA11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~27_cout ),
	.combout(),
	.cout(\LessThan0~29_cout ));
// synopsys translate_off
defparam \LessThan0~29 .lut_mask = 16'h002B;
defparam \LessThan0~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N30
cycloneive_lcell_comb \LessThan0~31 (
// Equation(s):
// \LessThan0~31_cout  = CARRY((\portA~27_combout  & ((!\LessThan0~29_cout ) # (!\portB~64_combout ))) # (!\portA~27_combout  & (!\portB~64_combout  & !\LessThan0~29_cout )))

	.dataa(portA10),
	.datab(portB16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~29_cout ),
	.combout(),
	.cout(\LessThan0~31_cout ));
// synopsys translate_off
defparam \LessThan0~31 .lut_mask = 16'h002B;
defparam \LessThan0~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N0
cycloneive_lcell_comb \LessThan0~33 (
// Equation(s):
// \LessThan0~33_cout  = CARRY((\portA~25_combout  & (\portB~62_combout  & !\LessThan0~31_cout )) # (!\portA~25_combout  & ((\portB~62_combout ) # (!\LessThan0~31_cout ))))

	.dataa(portA9),
	.datab(portB15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~31_cout ),
	.combout(),
	.cout(\LessThan0~33_cout ));
// synopsys translate_off
defparam \LessThan0~33 .lut_mask = 16'h004D;
defparam \LessThan0~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N2
cycloneive_lcell_comb \LessThan0~35 (
// Equation(s):
// \LessThan0~35_cout  = CARRY((\portB~59_combout  & (\portA~67_combout  & !\LessThan0~33_cout )) # (!\portB~59_combout  & ((\portA~67_combout ) # (!\LessThan0~33_cout ))))

	.dataa(portB14),
	.datab(portA31),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~33_cout ),
	.combout(),
	.cout(\LessThan0~35_cout ));
// synopsys translate_off
defparam \LessThan0~35 .lut_mask = 16'h004D;
defparam \LessThan0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N4
cycloneive_lcell_comb \LessThan0~37 (
// Equation(s):
// \LessThan0~37_cout  = CARRY((\portA~65_combout  & (\portB~56_combout  & !\LessThan0~35_cout )) # (!\portA~65_combout  & ((\portB~56_combout ) # (!\LessThan0~35_cout ))))

	.dataa(portA30),
	.datab(portB13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~35_cout ),
	.combout(),
	.cout(\LessThan0~37_cout ));
// synopsys translate_off
defparam \LessThan0~37 .lut_mask = 16'h004D;
defparam \LessThan0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N6
cycloneive_lcell_comb \LessThan0~39 (
// Equation(s):
// \LessThan0~39_cout  = CARRY((\portB~53_combout  & (\portA~63_combout  & !\LessThan0~37_cout )) # (!\portB~53_combout  & ((\portA~63_combout ) # (!\LessThan0~37_cout ))))

	.dataa(portB12),
	.datab(portA29),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~37_cout ),
	.combout(),
	.cout(\LessThan0~39_cout ));
// synopsys translate_off
defparam \LessThan0~39 .lut_mask = 16'h004D;
defparam \LessThan0~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N8
cycloneive_lcell_comb \LessThan0~41 (
// Equation(s):
// \LessThan0~41_cout  = CARRY((\portA~61_combout  & (\portB~50_combout  & !\LessThan0~39_cout )) # (!\portA~61_combout  & ((\portB~50_combout ) # (!\LessThan0~39_cout ))))

	.dataa(portA28),
	.datab(portB11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~39_cout ),
	.combout(),
	.cout(\LessThan0~41_cout ));
// synopsys translate_off
defparam \LessThan0~41 .lut_mask = 16'h004D;
defparam \LessThan0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N10
cycloneive_lcell_comb \LessThan0~43 (
// Equation(s):
// \LessThan0~43_cout  = CARRY((\portB~47_combout  & (\portA~59_combout  & !\LessThan0~41_cout )) # (!\portB~47_combout  & ((\portA~59_combout ) # (!\LessThan0~41_cout ))))

	.dataa(portB10),
	.datab(portA27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~41_cout ),
	.combout(),
	.cout(\LessThan0~43_cout ));
// synopsys translate_off
defparam \LessThan0~43 .lut_mask = 16'h004D;
defparam \LessThan0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N12
cycloneive_lcell_comb \LessThan0~45 (
// Equation(s):
// \LessThan0~45_cout  = CARRY((\portA~57_combout  & (\portB~44_combout  & !\LessThan0~43_cout )) # (!\portA~57_combout  & ((\portB~44_combout ) # (!\LessThan0~43_cout ))))

	.dataa(portA26),
	.datab(portB9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~43_cout ),
	.combout(),
	.cout(\LessThan0~45_cout ));
// synopsys translate_off
defparam \LessThan0~45 .lut_mask = 16'h004D;
defparam \LessThan0~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N14
cycloneive_lcell_comb \LessThan0~47 (
// Equation(s):
// \LessThan0~47_cout  = CARRY((\portA~55_combout  & ((!\LessThan0~45_cout ) # (!\portB~41_combout ))) # (!\portA~55_combout  & (!\portB~41_combout  & !\LessThan0~45_cout )))

	.dataa(portA25),
	.datab(portB8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~45_cout ),
	.combout(),
	.cout(\LessThan0~47_cout ));
// synopsys translate_off
defparam \LessThan0~47 .lut_mask = 16'h002B;
defparam \LessThan0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N16
cycloneive_lcell_comb \LessThan0~49 (
// Equation(s):
// \LessThan0~49_cout  = CARRY((\portB~38_combout  & ((!\LessThan0~47_cout ) # (!\portA~53_combout ))) # (!\portB~38_combout  & (!\portA~53_combout  & !\LessThan0~47_cout )))

	.dataa(portB7),
	.datab(portA24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~47_cout ),
	.combout(),
	.cout(\LessThan0~49_cout ));
// synopsys translate_off
defparam \LessThan0~49 .lut_mask = 16'h002B;
defparam \LessThan0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N18
cycloneive_lcell_comb \LessThan0~51 (
// Equation(s):
// \LessThan0~51_cout  = CARRY((\portB~35_combout  & (\portA~51_combout  & !\LessThan0~49_cout )) # (!\portB~35_combout  & ((\portA~51_combout ) # (!\LessThan0~49_cout ))))

	.dataa(portB6),
	.datab(portA23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~49_cout ),
	.combout(),
	.cout(\LessThan0~51_cout ));
// synopsys translate_off
defparam \LessThan0~51 .lut_mask = 16'h004D;
defparam \LessThan0~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N20
cycloneive_lcell_comb \LessThan0~53 (
// Equation(s):
// \LessThan0~53_cout  = CARRY((\portA~49_combout  & (\portB~32_combout  & !\LessThan0~51_cout )) # (!\portA~49_combout  & ((\portB~32_combout ) # (!\LessThan0~51_cout ))))

	.dataa(portA22),
	.datab(portB5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~51_cout ),
	.combout(),
	.cout(\LessThan0~53_cout ));
// synopsys translate_off
defparam \LessThan0~53 .lut_mask = 16'h004D;
defparam \LessThan0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N22
cycloneive_lcell_comb \LessThan0~55 (
// Equation(s):
// \LessThan0~55_cout  = CARRY((\portA~47_combout  & ((!\LessThan0~53_cout ) # (!\portB~29_combout ))) # (!\portA~47_combout  & (!\portB~29_combout  & !\LessThan0~53_cout )))

	.dataa(portA21),
	.datab(portB4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~53_cout ),
	.combout(),
	.cout(\LessThan0~55_cout ));
// synopsys translate_off
defparam \LessThan0~55 .lut_mask = 16'h002B;
defparam \LessThan0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N24
cycloneive_lcell_comb \LessThan0~57 (
// Equation(s):
// \LessThan0~57_cout  = CARRY((\portA~45_combout  & (\portB~26_combout  & !\LessThan0~55_cout )) # (!\portA~45_combout  & ((\portB~26_combout ) # (!\LessThan0~55_cout ))))

	.dataa(portA20),
	.datab(portB3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~55_cout ),
	.combout(),
	.cout(\LessThan0~57_cout ));
// synopsys translate_off
defparam \LessThan0~57 .lut_mask = 16'h004D;
defparam \LessThan0~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N26
cycloneive_lcell_comb \LessThan0~59 (
// Equation(s):
// \LessThan0~59_cout  = CARRY((\portA~41_combout  & ((!\LessThan0~57_cout ) # (!\portB~23_combout ))) # (!\portA~41_combout  & (!\portB~23_combout  & !\LessThan0~57_cout )))

	.dataa(portA18),
	.datab(portB2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~57_cout ),
	.combout(),
	.cout(\LessThan0~59_cout ));
// synopsys translate_off
defparam \LessThan0~59 .lut_mask = 16'h002B;
defparam \LessThan0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N28
cycloneive_lcell_comb \LessThan0~61 (
// Equation(s):
// \LessThan0~61_cout  = CARRY((\portB~20_combout  & ((!\LessThan0~59_cout ) # (!\portA~43_combout ))) # (!\portB~20_combout  & (!\portA~43_combout  & !\LessThan0~59_cout )))

	.dataa(portB1),
	.datab(portA19),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~59_cout ),
	.combout(),
	.cout(\LessThan0~61_cout ));
// synopsys translate_off
defparam \LessThan0~61 .lut_mask = 16'h002B;
defparam \LessThan0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N30
cycloneive_lcell_comb \LessThan0~62 (
// Equation(s):
// \LessThan0~62_combout  = (\portB~17_combout  & (\LessThan0~61_cout  & \portA~39_combout )) # (!\portB~17_combout  & ((\LessThan0~61_cout ) # (\portA~39_combout )))

	.dataa(gnd),
	.datab(portB),
	.datac(gnd),
	.datad(portA17),
	.cin(\LessThan0~61_cout ),
	.combout(\LessThan0~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan0~62 .lut_mask = 16'hF330;
defparam \LessThan0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N18
cycloneive_lcell_comb \Selector31~1 (
// Equation(s):
// \Selector31~1_combout  = (ALUOp_EX[1] & ((ALUOp_EX[0] & (\LessThan1~62_combout )) # (!ALUOp_EX[0] & ((\LessThan0~62_combout )))))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_1),
	.datac(\LessThan1~62_combout ),
	.datad(\LessThan0~62_combout ),
	.cin(gnd),
	.combout(\Selector31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~1 .lut_mask = 16'hC480;
defparam \Selector31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N24
cycloneive_lcell_comb \ShiftRight0~40 (
// Equation(s):
// \ShiftRight0~40_combout  = (\portB~92_combout  & ((\portA~35_combout ))) # (!\portB~92_combout  & (\portA~36_combout ))

	.dataa(gnd),
	.datab(portA15),
	.datac(portA14),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~40 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N10
cycloneive_lcell_comb \ShiftRight0~41 (
// Equation(s):
// \ShiftRight0~41_combout  = (\portB~92_combout  & ((\portA~37_combout ))) # (!\portB~92_combout  & (\portA~17_combout ))

	.dataa(gnd),
	.datab(portA5),
	.datac(portA16),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~41 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N16
cycloneive_lcell_comb \ShiftRight0~42 (
// Equation(s):
// \ShiftRight0~42_combout  = (\portB~97_combout  & (\ShiftRight0~40_combout )) # (!\portB~97_combout  & ((\ShiftRight0~41_combout )))

	.dataa(portB30),
	.datab(\ShiftRight0~40_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~41_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~42 .lut_mask = 16'hDD88;
defparam \ShiftRight0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N6
cycloneive_lcell_comb \ShiftRight0~38 (
// Equation(s):
// \ShiftRight0~38_combout  = (\portB~92_combout  & (\portA~31_combout )) # (!\portB~92_combout  & ((\portA~33_combout )))

	.dataa(gnd),
	.datab(portA12),
	.datac(portA13),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~38 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N28
cycloneive_lcell_comb \ShiftRight0~37 (
// Equation(s):
// \ShiftRight0~37_combout  = (\portB~92_combout  & (\portA~27_combout )) # (!\portB~92_combout  & ((\portA~29_combout )))

	.dataa(portA10),
	.datab(gnd),
	.datac(portB29),
	.datad(portA11),
	.cin(gnd),
	.combout(\ShiftRight0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~37 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N20
cycloneive_lcell_comb \ShiftRight0~39 (
// Equation(s):
// \ShiftRight0~39_combout  = (\portB~97_combout  & ((\ShiftRight0~37_combout ))) # (!\portB~97_combout  & (\ShiftRight0~38_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftRight0~38_combout ),
	.datad(\ShiftRight0~37_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~39 .lut_mask = 16'hFA50;
defparam \ShiftRight0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N12
cycloneive_lcell_comb \ShiftRight0~43 (
// Equation(s):
// \ShiftRight0~43_combout  = (\portB~100_combout  & ((\ShiftRight0~39_combout ))) # (!\portB~100_combout  & (\ShiftRight0~42_combout ))

	.dataa(portB31),
	.datab(gnd),
	.datac(\ShiftRight0~42_combout ),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~43 .lut_mask = 16'hFA50;
defparam \ShiftRight0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N30
cycloneive_lcell_comb \ShiftRight0~31 (
// Equation(s):
// \ShiftRight0~31_combout  = (\portB~92_combout  & (\portA~16_combout )) # (!\portB~92_combout  & ((\portA~9_combout )))

	.dataa(gnd),
	.datab(portA4),
	.datac(portB29),
	.datad(portA),
	.cin(gnd),
	.combout(\ShiftRight0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~31 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N2
cycloneive_lcell_comb \ShiftRight0~30 (
// Equation(s):
// \ShiftRight0~30_combout  = (!\portB~97_combout  & ((\portB~92_combout  & (\portA~12_combout )) # (!\portB~92_combout  & ((\portA~69_combout )))))

	.dataa(portA1),
	.datab(portB30),
	.datac(portA32),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~30 .lut_mask = 16'h2230;
defparam \ShiftRight0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N16
cycloneive_lcell_comb \ShiftRight0~32 (
// Equation(s):
// \ShiftRight0~32_combout  = (!\portB~100_combout  & ((\ShiftRight0~30_combout ) # ((\portB~97_combout  & \ShiftRight0~31_combout ))))

	.dataa(portB31),
	.datab(portB30),
	.datac(\ShiftRight0~31_combout ),
	.datad(\ShiftRight0~30_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~32 .lut_mask = 16'h5540;
defparam \ShiftRight0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N6
cycloneive_lcell_comb \ShiftRight0~36 (
// Equation(s):
// \ShiftRight0~36_combout  = (!\portB~103_combout  & ((\ShiftRight0~32_combout ) # ((\ShiftRight0~35_combout  & \portB~100_combout ))))

	.dataa(\ShiftRight0~35_combout ),
	.datab(\ShiftRight0~32_combout ),
	.datac(portB32),
	.datad(portB31),
	.cin(gnd),
	.combout(\ShiftRight0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~36 .lut_mask = 16'h0E0C;
defparam \ShiftRight0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N26
cycloneive_lcell_comb \ShiftRight0~44 (
// Equation(s):
// \ShiftRight0~44_combout  = (!\portB~107_combout  & ((\ShiftRight0~36_combout ) # ((\portB~103_combout  & \ShiftRight0~43_combout ))))

	.dataa(portB33),
	.datab(portB32),
	.datac(\ShiftRight0~43_combout ),
	.datad(\ShiftRight0~36_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~44 .lut_mask = 16'h5540;
defparam \ShiftRight0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N16
cycloneive_lcell_comb \ShiftRight0~53 (
// Equation(s):
// \ShiftRight0~53_combout  = (\portB~92_combout  & ((\portA~59_combout ))) # (!\portB~92_combout  & (\portA~61_combout ))

	.dataa(gnd),
	.datab(portA28),
	.datac(portA27),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~53 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N30
cycloneive_lcell_comb \ShiftRight0~52 (
// Equation(s):
// \ShiftRight0~52_combout  = (\portB~92_combout  & (\portA~55_combout )) # (!\portB~92_combout  & ((\portA~57_combout )))

	.dataa(gnd),
	.datab(portA25),
	.datac(portB29),
	.datad(portA26),
	.cin(gnd),
	.combout(\ShiftRight0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~52 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N18
cycloneive_lcell_comb \ShiftRight0~54 (
// Equation(s):
// \ShiftRight0~54_combout  = (\portB~97_combout  & ((\ShiftRight0~52_combout ))) # (!\portB~97_combout  & (\ShiftRight0~53_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~53_combout ),
	.datac(portB30),
	.datad(\ShiftRight0~52_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~54 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N28
cycloneive_lcell_comb \Selector23~0 (
// Equation(s):
// \Selector23~0_combout  = (\portB~100_combout  & ((\ShiftRight0~54_combout ))) # (!\portB~100_combout  & (\ShiftRight0~57_combout ))

	.dataa(\ShiftRight0~57_combout ),
	.datab(\ShiftRight0~54_combout ),
	.datac(gnd),
	.datad(portB31),
	.cin(gnd),
	.combout(\Selector23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~0 .lut_mask = 16'hCCAA;
defparam \Selector23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N0
cycloneive_lcell_comb \ShiftRight0~48 (
// Equation(s):
// \ShiftRight0~48_combout  = (\portB~92_combout  & (\portA~47_combout )) # (!\portB~92_combout  & ((\portA~49_combout )))

	.dataa(portA21),
	.datab(gnd),
	.datac(portB29),
	.datad(portA22),
	.cin(gnd),
	.combout(\ShiftRight0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~48 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N2
cycloneive_lcell_comb \ShiftRight0~49 (
// Equation(s):
// \ShiftRight0~49_combout  = (\portB~92_combout  & ((\portA~51_combout ))) # (!\portB~92_combout  & (\portA~53_combout ))

	.dataa(gnd),
	.datab(portA24),
	.datac(portA23),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~49 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N8
cycloneive_lcell_comb \ShiftRight0~50 (
// Equation(s):
// \ShiftRight0~50_combout  = (\portB~97_combout  & (\ShiftRight0~48_combout )) # (!\portB~97_combout  & ((\ShiftRight0~49_combout )))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftRight0~48_combout ),
	.datad(\ShiftRight0~49_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~50 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N8
cycloneive_lcell_comb \ShiftRight0~46 (
// Equation(s):
// \ShiftRight0~46_combout  = (\portB~92_combout  & (\portA~41_combout )) # (!\portB~92_combout  & ((\portA~45_combout )))

	.dataa(portA18),
	.datab(portB29),
	.datac(gnd),
	.datad(portA20),
	.cin(gnd),
	.combout(\ShiftRight0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~46 .lut_mask = 16'hBB88;
defparam \ShiftRight0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N10
cycloneive_lcell_comb \ShiftRight0~45 (
// Equation(s):
// \ShiftRight0~45_combout  = (\portB~92_combout  & ((\portA~39_combout ))) # (!\portB~92_combout  & (\portA~43_combout ))

	.dataa(portA19),
	.datab(portB29),
	.datac(portA17),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~45 .lut_mask = 16'hE2E2;
defparam \ShiftRight0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N22
cycloneive_lcell_comb \ShiftRight0~47 (
// Equation(s):
// \ShiftRight0~47_combout  = (\portB~97_combout  & ((\ShiftRight0~45_combout ))) # (!\portB~97_combout  & (\ShiftRight0~46_combout ))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftRight0~46_combout ),
	.datad(\ShiftRight0~45_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~47 .lut_mask = 16'hFC30;
defparam \ShiftRight0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N14
cycloneive_lcell_comb \ShiftRight0~51 (
// Equation(s):
// \ShiftRight0~51_combout  = (\portB~100_combout  & ((\ShiftRight0~47_combout ))) # (!\portB~100_combout  & (\ShiftRight0~50_combout ))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftRight0~50_combout ),
	.datad(\ShiftRight0~47_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~51 .lut_mask = 16'hFC30;
defparam \ShiftRight0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N24
cycloneive_lcell_comb \ShiftRight0~58 (
// Equation(s):
// \ShiftRight0~58_combout  = (\portB~103_combout  & ((\ShiftRight0~51_combout ))) # (!\portB~103_combout  & (\Selector23~0_combout ))

	.dataa(gnd),
	.datab(portB32),
	.datac(\Selector23~0_combout ),
	.datad(\ShiftRight0~51_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~58 .lut_mask = 16'hFC30;
defparam \ShiftRight0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N30
cycloneive_lcell_comb \ShiftLeft0~15 (
// Equation(s):
// \ShiftLeft0~15_combout  = (\portB~100_combout ) # ((\portB~97_combout ) # ((\portB~103_combout ) # (\portB~92_combout )))

	.dataa(portB31),
	.datab(portB30),
	.datac(portB32),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~15 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N10
cycloneive_lcell_comb \Selector31~7 (
// Equation(s):
// \Selector31~7_combout  = (\Selector0~2_combout ) # ((\Selector0~3_combout  & \portB~92_combout ))

	.dataa(\Selector0~2_combout ),
	.datab(\Selector0~3_combout ),
	.datac(gnd),
	.datad(portB29),
	.cin(gnd),
	.combout(\Selector31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~7 .lut_mask = 16'hEEAA;
defparam \Selector31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N26
cycloneive_lcell_comb \Selector0~10 (
// Equation(s):
// \Selector0~10_combout  = (!ALUOp_EX[0] & (ALUOp_EX[2] & (!ALUOp_EX[3] & ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~10 .lut_mask = 16'h0400;
defparam \Selector0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N10
cycloneive_lcell_comb \Selector0~8 (
// Equation(s):
// \Selector0~8_combout  = (!ALUOp_EX[3] & (ALUOp_EX[2] & (ALUOp_EX[0] & !ALUOp_EX[1])))

	.dataa(ALUOp_EX_3),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_0),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~8 .lut_mask = 16'h0040;
defparam \Selector0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N24
cycloneive_lcell_comb \Selector28~4 (
// Equation(s):
// \Selector28~4_combout  = (\portA~16_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \portB~103_combout ))))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector0~8_combout ),
	.datac(portB32),
	.datad(portA4),
	.cin(gnd),
	.combout(\Selector28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~4 .lut_mask = 16'hEC00;
defparam \Selector28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N26
cycloneive_lcell_comb \Selector28~5 (
// Equation(s):
// \Selector28~5_combout  = (\Selector28~4_combout ) # ((\Selector0~10_combout  & (\portB~103_combout  $ (\portA~16_combout ))))

	.dataa(portB32),
	.datab(portA4),
	.datac(\Selector0~10_combout ),
	.datad(\Selector28~4_combout ),
	.cin(gnd),
	.combout(\Selector28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~5 .lut_mask = 16'hFF60;
defparam \Selector28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N26
cycloneive_lcell_comb \ShiftLeft0~17 (
// Equation(s):
// \ShiftLeft0~17_combout  = (!\portB~100_combout  & !\portB~103_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(portB31),
	.datad(portB32),
	.cin(gnd),
	.combout(\ShiftLeft0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~17 .lut_mask = 16'h000F;
defparam \ShiftLeft0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N2
cycloneive_lcell_comb \ShiftLeft0~16 (
// Equation(s):
// \ShiftLeft0~16_combout  = (\ShiftLeft0~7_combout ) # ((\ShiftLeft0~6_combout ) # (\ShiftLeft0~10_combout ))

	.dataa(\ShiftLeft0~7_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~6_combout ),
	.datad(\ShiftLeft0~10_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~16 .lut_mask = 16'hFFFA;
defparam \ShiftLeft0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N20
cycloneive_lcell_comb \Selector29~0 (
// Equation(s):
// \Selector29~0_combout  = (\Selector0~14_combout  & (!\portB~107_combout  & (\ShiftLeft0~17_combout  & !\ShiftLeft0~16_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(portB33),
	.datac(\ShiftLeft0~17_combout ),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~0 .lut_mask = 16'h0020;
defparam \Selector29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N8
cycloneive_lcell_comb \ShiftLeft0~18 (
// Equation(s):
// \ShiftLeft0~18_combout  = (\portB~92_combout  & ((\portA~9_combout ))) # (!\portB~92_combout  & (\portA~16_combout ))

	.dataa(gnd),
	.datab(portA4),
	.datac(portB29),
	.datad(portA),
	.cin(gnd),
	.combout(\ShiftLeft0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~18 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N26
cycloneive_lcell_comb \ShiftLeft0~19 (
// Equation(s):
// \ShiftLeft0~19_combout  = (\portB~97_combout  & ((\ShiftLeft0~13_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~18_combout ))

	.dataa(portB30),
	.datab(\ShiftLeft0~18_combout ),
	.datac(\ShiftLeft0~13_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~19 .lut_mask = 16'hE4E4;
defparam \ShiftLeft0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N28
cycloneive_lcell_comb \Selector0~13 (
// Equation(s):
// \Selector0~13_combout  = (!ALUOp_EX[3] & (ALUOp_EX[2] & (ALUOp_EX[0] & ALUOp_EX[1])))

	.dataa(ALUOp_EX_3),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_0),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~13 .lut_mask = 16'h4000;
defparam \Selector0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N20
cycloneive_lcell_comb \Selector28~7 (
// Equation(s):
// \Selector28~7_combout  = (\Selector0~13_combout  & ((fuifforward_A_11 & (!\wdat_WB[3]~65_combout )) # (!fuifforward_A_11 & ((!\portA~15_combout )))))

	.dataa(wdat_WB_3),
	.datab(portA3),
	.datac(\Selector0~13_combout ),
	.datad(fuifforward_A_1),
	.cin(gnd),
	.combout(\Selector28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~7 .lut_mask = 16'h5030;
defparam \Selector28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N6
cycloneive_lcell_comb \Selector0~11 (
// Equation(s):
// \Selector0~11_combout  = (!ALUOp_EX[2] & (ALUOp_EX[0] & (ALUOp_EX[1] & !ALUOp_EX[3])))

	.dataa(ALUOp_EX_2),
	.datab(ALUOp_EX_0),
	.datac(ALUOp_EX_1),
	.datad(ALUOp_EX_3),
	.cin(gnd),
	.combout(\Selector0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~11 .lut_mask = 16'h0040;
defparam \Selector0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N4
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = ((\portB~100_combout  $ (\portA~9_combout  $ (!\Add0~3 )))) # (GND)
// \Add0~5  = CARRY((\portB~100_combout  & ((\portA~9_combout ) # (!\Add0~3 ))) # (!\portB~100_combout  & (\portA~9_combout  & !\Add0~3 )))

	.dataa(portB31),
	.datab(portA),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'h698E;
defparam \Add0~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N6
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = (\portA~16_combout  & ((\portB~103_combout  & (\Add0~5  & VCC)) # (!\portB~103_combout  & (!\Add0~5 )))) # (!\portA~16_combout  & ((\portB~103_combout  & (!\Add0~5 )) # (!\portB~103_combout  & ((\Add0~5 ) # (GND)))))
// \Add0~7  = CARRY((\portA~16_combout  & (!\portB~103_combout  & !\Add0~5 )) # (!\portA~16_combout  & ((!\Add0~5 ) # (!\portB~103_combout ))))

	.dataa(portA4),
	.datab(portB32),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h9617;
defparam \Add0~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N4
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((\portB~100_combout  $ (\portA~9_combout  $ (\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((\portB~100_combout  & (\portA~9_combout  & !\Add1~3 )) # (!\portB~100_combout  & ((\portA~9_combout ) # (!\Add1~3 ))))

	.dataa(portB31),
	.datab(portA),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h964D;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N6
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (\portA~16_combout  & ((\portB~103_combout  & (!\Add1~5 )) # (!\portB~103_combout  & (\Add1~5  & VCC)))) # (!\portA~16_combout  & ((\portB~103_combout  & ((\Add1~5 ) # (GND))) # (!\portB~103_combout  & (!\Add1~5 ))))
// \Add1~7  = CARRY((\portA~16_combout  & (\portB~103_combout  & !\Add1~5 )) # (!\portA~16_combout  & ((\portB~103_combout ) # (!\Add1~5 ))))

	.dataa(portA4),
	.datab(portB32),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h694D;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N28
cycloneive_lcell_comb \Selector28~6 (
// Equation(s):
// \Selector28~6_combout  = (\Selector0~12_combout  & ((\Add0~6_combout ) # ((\Selector0~11_combout  & \Add1~6_combout )))) # (!\Selector0~12_combout  & (\Selector0~11_combout  & ((\Add1~6_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Add0~6_combout ),
	.datad(\Add1~6_combout ),
	.cin(gnd),
	.combout(\Selector28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~6 .lut_mask = 16'hECA0;
defparam \Selector28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N10
cycloneive_lcell_comb \Selector28~8 (
// Equation(s):
// \Selector28~8_combout  = (\Selector28~6_combout ) # ((\portB~103_combout  & (\Selector0~8_combout )) # (!\portB~103_combout  & ((\Selector28~7_combout ))))

	.dataa(portB32),
	.datab(\Selector0~8_combout ),
	.datac(\Selector28~7_combout ),
	.datad(\Selector28~6_combout ),
	.cin(gnd),
	.combout(\Selector28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~8 .lut_mask = 16'hFFD8;
defparam \Selector28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N22
cycloneive_lcell_comb \Selector28~9 (
// Equation(s):
// \Selector28~9_combout  = (\Selector28~5_combout ) # ((\Selector28~8_combout ) # ((\Selector29~0_combout  & \ShiftLeft0~19_combout )))

	.dataa(\Selector28~5_combout ),
	.datab(\Selector29~0_combout ),
	.datac(\ShiftLeft0~19_combout ),
	.datad(\Selector28~8_combout ),
	.cin(gnd),
	.combout(\Selector28~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~9 .lut_mask = 16'hFFEA;
defparam \Selector28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N14
cycloneive_lcell_comb \Selector12~4 (
// Equation(s):
// \Selector12~4_combout  = (!ALUOp_EX[2] & !ALUOp_EX[3])

	.dataa(gnd),
	.datab(ALUOp_EX_2),
	.datac(gnd),
	.datad(ALUOp_EX_3),
	.cin(gnd),
	.combout(\Selector12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~4 .lut_mask = 16'h0033;
defparam \Selector12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N16
cycloneive_lcell_comb \Selector12~5 (
// Equation(s):
// \Selector12~5_combout  = (!ALUOp_EX[1] & (\Selector12~4_combout  & (!\ShiftLeft0~12_combout  & !\ShiftLeft0~6_combout )))

	.dataa(ALUOp_EX_1),
	.datab(\Selector12~4_combout ),
	.datac(\ShiftLeft0~12_combout ),
	.datad(\ShiftLeft0~6_combout ),
	.cin(gnd),
	.combout(\Selector12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~5 .lut_mask = 16'h0004;
defparam \Selector12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N24
cycloneive_lcell_comb \Selector16~0 (
// Equation(s):
// \Selector16~0_combout  = (\portB~107_combout  & (ALUOp_EX[0] & \Selector12~5_combout ))

	.dataa(gnd),
	.datab(portB33),
	.datac(ALUOp_EX_0),
	.datad(\Selector12~5_combout ),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~0 .lut_mask = 16'hC000;
defparam \Selector16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N4
cycloneive_lcell_comb \ShiftRight0~67 (
// Equation(s):
// \ShiftRight0~67_combout  = (\portB~97_combout  & ((\ShiftRight0~20_combout ))) # (!\portB~97_combout  & (\ShiftRight0~23_combout ))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftRight0~23_combout ),
	.datad(\ShiftRight0~20_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~67 .lut_mask = 16'hFC30;
defparam \ShiftRight0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N8
cycloneive_lcell_comb \ShiftRight0~68 (
// Equation(s):
// \ShiftRight0~68_combout  = (\portB~97_combout  & (\ShiftRight0~24_combout )) # (!\portB~97_combout  & ((\ShiftRight0~26_combout )))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftRight0~24_combout ),
	.datad(\ShiftRight0~26_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~68 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N14
cycloneive_lcell_comb \Selector20~0 (
// Equation(s):
// \Selector20~0_combout  = (\portB~100_combout  & (\ShiftRight0~67_combout )) # (!\portB~100_combout  & ((\ShiftRight0~68_combout )))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftRight0~67_combout ),
	.datad(\ShiftRight0~68_combout ),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~0 .lut_mask = 16'hF3C0;
defparam \Selector20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N22
cycloneive_lcell_comb \ShiftRight0~63 (
// Equation(s):
// \ShiftRight0~63_combout  = (\portA~39_combout  & (!\portB~97_combout  & !\portB~92_combout ))

	.dataa(portA17),
	.datab(gnd),
	.datac(portB30),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~63 .lut_mask = 16'h000A;
defparam \ShiftRight0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N8
cycloneive_lcell_comb \ShiftRight0~64 (
// Equation(s):
// \ShiftRight0~64_combout  = (\portB~97_combout  & ((\portB~92_combout  & ((\portA~43_combout ))) # (!\portB~92_combout  & (\portA~41_combout ))))

	.dataa(portA18),
	.datab(portA19),
	.datac(portB30),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~64 .lut_mask = 16'hC0A0;
defparam \ShiftRight0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N10
cycloneive_lcell_comb \ShiftRight0~65 (
// Equation(s):
// \ShiftRight0~65_combout  = (\ShiftRight0~64_combout ) # ((!\portB~97_combout  & \ShiftRight0~19_combout ))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftRight0~64_combout ),
	.datad(\ShiftRight0~19_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~65 .lut_mask = 16'hF3F0;
defparam \ShiftRight0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N4
cycloneive_lcell_comb \ShiftRight0~66 (
// Equation(s):
// \ShiftRight0~66_combout  = (\portB~100_combout  & (\ShiftRight0~63_combout )) # (!\portB~100_combout  & ((\ShiftRight0~65_combout )))

	.dataa(portB31),
	.datab(gnd),
	.datac(\ShiftRight0~63_combout ),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~66 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N24
cycloneive_lcell_comb \ShiftRight0~69 (
// Equation(s):
// \ShiftRight0~69_combout  = (\portB~103_combout  & ((\ShiftRight0~66_combout ))) # (!\portB~103_combout  & (\Selector20~0_combout ))

	.dataa(gnd),
	.datab(portB32),
	.datac(\Selector20~0_combout ),
	.datad(\ShiftRight0~66_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~69 .lut_mask = 16'hFC30;
defparam \ShiftRight0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N14
cycloneive_lcell_comb \Selector12~19 (
// Equation(s):
// \Selector12~19_combout  = (!ALUOp_EX[2] & (!\ShiftLeft0~6_combout  & (!\ShiftLeft0~12_combout  & !ALUOp_EX[3])))

	.dataa(ALUOp_EX_2),
	.datab(\ShiftLeft0~6_combout ),
	.datac(\ShiftLeft0~12_combout ),
	.datad(ALUOp_EX_3),
	.cin(gnd),
	.combout(\Selector12~19_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~19 .lut_mask = 16'h0001;
defparam \Selector12~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N16
cycloneive_lcell_comb \Selector28~0 (
// Equation(s):
// \Selector28~0_combout  = (ALUOp_EX[0] & (!ALUOp_EX[1] & ((\ShiftLeft0~16_combout ) # (!\portB~107_combout ))))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_1),
	.datac(portB33),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~0 .lut_mask = 16'h2202;
defparam \Selector28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N30
cycloneive_lcell_comb \ShiftRight0~59 (
// Equation(s):
// \ShiftRight0~59_combout  = (\portB~97_combout  & ((\ShiftRight0~13_combout ))) # (!\portB~97_combout  & (\ShiftRight0~5_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftRight0~5_combout ),
	.datad(\ShiftRight0~13_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~59 .lut_mask = 16'hFA50;
defparam \ShiftRight0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N8
cycloneive_lcell_comb \Selector2~2 (
// Equation(s):
// \Selector2~2_combout  = (\portB~103_combout ) # ((!\portB~100_combout  & \portB~97_combout ))

	.dataa(gnd),
	.datab(portB32),
	.datac(portB31),
	.datad(portB30),
	.cin(gnd),
	.combout(\Selector2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~2 .lut_mask = 16'hCFCC;
defparam \Selector2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N0
cycloneive_lcell_comb \Selector28~1 (
// Equation(s):
// \Selector28~1_combout  = (\ShiftLeft0~17_combout  & (\ShiftRight0~3_combout  & ((!\Selector2~2_combout )))) # (!\ShiftLeft0~17_combout  & (((\ShiftRight0~59_combout ) # (\Selector2~2_combout ))))

	.dataa(\ShiftLeft0~17_combout ),
	.datab(\ShiftRight0~3_combout ),
	.datac(\ShiftRight0~59_combout ),
	.datad(\Selector2~2_combout ),
	.cin(gnd),
	.combout(\Selector28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~1 .lut_mask = 16'h55D8;
defparam \Selector28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N8
cycloneive_lcell_comb \ShiftRight0~9 (
// Equation(s):
// \ShiftRight0~9_combout  = (\portB~92_combout  & (\portA~25_combout )) # (!\portB~92_combout  & ((\portA~27_combout )))

	.dataa(gnd),
	.datab(portA9),
	.datac(portA10),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~9 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N30
cycloneive_lcell_comb \ShiftRight0~60 (
// Equation(s):
// \ShiftRight0~60_combout  = (\portB~97_combout  & (\ShiftRight0~27_combout )) # (!\portB~97_combout  & ((\ShiftRight0~9_combout )))

	.dataa(\ShiftRight0~27_combout ),
	.datab(gnd),
	.datac(portB30),
	.datad(\ShiftRight0~9_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~60 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N30
cycloneive_lcell_comb \ShiftRight0~10 (
// Equation(s):
// \ShiftRight0~10_combout  = (\portB~92_combout  & ((\portA~29_combout ))) # (!\portB~92_combout  & (\portA~31_combout ))

	.dataa(gnd),
	.datab(portA12),
	.datac(portA11),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~10 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N10
cycloneive_lcell_comb \ShiftRight0~61 (
// Equation(s):
// \ShiftRight0~61_combout  = (\portB~97_combout  & ((\ShiftRight0~10_combout ))) # (!\portB~97_combout  & (\ShiftRight0~12_combout ))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftRight0~12_combout ),
	.datad(\ShiftRight0~10_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~61 .lut_mask = 16'hFC30;
defparam \ShiftRight0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N16
cycloneive_lcell_comb \ShiftRight0~62 (
// Equation(s):
// \ShiftRight0~62_combout  = (\portB~100_combout  & (\ShiftRight0~60_combout )) # (!\portB~100_combout  & ((\ShiftRight0~61_combout )))

	.dataa(portB31),
	.datab(gnd),
	.datac(\ShiftRight0~60_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~62 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N4
cycloneive_lcell_comb \Selector28~2 (
// Equation(s):
// \Selector28~2_combout  = (\Selector2~2_combout  & ((\Selector28~1_combout  & ((\ShiftRight0~62_combout ))) # (!\Selector28~1_combout  & (\ShiftRight0~6_combout )))) # (!\Selector2~2_combout  & (((\Selector28~1_combout ))))

	.dataa(\Selector2~2_combout ),
	.datab(\ShiftRight0~6_combout ),
	.datac(\Selector28~1_combout ),
	.datad(\ShiftRight0~62_combout ),
	.cin(gnd),
	.combout(\Selector28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~2 .lut_mask = 16'hF858;
defparam \Selector28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N2
cycloneive_lcell_comb \Selector28~3 (
// Equation(s):
// \Selector28~3_combout  = (\Selector12~19_combout  & (\Selector28~0_combout  & \Selector28~2_combout ))

	.dataa(\Selector12~19_combout ),
	.datab(\Selector28~0_combout ),
	.datac(gnd),
	.datad(\Selector28~2_combout ),
	.cin(gnd),
	.combout(\Selector28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~3 .lut_mask = 16'h8800;
defparam \Selector28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N18
cycloneive_lcell_comb \ShiftRight0~34 (
// Equation(s):
// \ShiftRight0~34_combout  = (\portB~92_combout  & ((\portA~23_combout ))) # (!\portB~92_combout  & (\portA~14_combout ))

	.dataa(gnd),
	.datab(portA2),
	.datac(portB29),
	.datad(portA8),
	.cin(gnd),
	.combout(\ShiftRight0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~34 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N22
cycloneive_lcell_comb \ShiftRight0~72 (
// Equation(s):
// \ShiftRight0~72_combout  = (\portB~97_combout  & (\ShiftRight0~38_combout )) # (!\portB~97_combout  & ((\ShiftRight0~40_combout )))

	.dataa(\ShiftRight0~38_combout ),
	.datab(gnd),
	.datac(portB30),
	.datad(\ShiftRight0~40_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~72 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N24
cycloneive_lcell_comb \ShiftRight0~71 (
// Equation(s):
// \ShiftRight0~71_combout  = (\portB~97_combout  & (\ShiftRight0~56_combout )) # (!\portB~97_combout  & ((\ShiftRight0~37_combout )))

	.dataa(\ShiftRight0~56_combout ),
	.datab(\ShiftRight0~37_combout ),
	.datac(gnd),
	.datad(portB30),
	.cin(gnd),
	.combout(\ShiftRight0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~71 .lut_mask = 16'hAACC;
defparam \ShiftRight0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N0
cycloneive_lcell_comb \ShiftRight0~73 (
// Equation(s):
// \ShiftRight0~73_combout  = (\portB~100_combout  & ((\ShiftRight0~71_combout ))) # (!\portB~100_combout  & (\ShiftRight0~72_combout ))

	.dataa(portB31),
	.datab(gnd),
	.datac(\ShiftRight0~72_combout ),
	.datad(\ShiftRight0~71_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~73 .lut_mask = 16'hFA50;
defparam \ShiftRight0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N14
cycloneive_lcell_comb \Selector29~2 (
// Equation(s):
// \Selector29~2_combout  = (\Selector29~1_combout  & (((\ShiftRight0~73_combout )) # (!\Selector2~2_combout ))) # (!\Selector29~1_combout  & (\Selector2~2_combout  & (\ShiftRight0~34_combout )))

	.dataa(\Selector29~1_combout ),
	.datab(\Selector2~2_combout ),
	.datac(\ShiftRight0~34_combout ),
	.datad(\ShiftRight0~73_combout ),
	.cin(gnd),
	.combout(\Selector29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~2 .lut_mask = 16'hEA62;
defparam \Selector29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N8
cycloneive_lcell_comb \Selector29~3 (
// Equation(s):
// \Selector29~3_combout  = (\Selector12~4_combout  & (\Selector29~2_combout  & (!\ShiftLeft0~16_combout  & \Selector28~0_combout )))

	.dataa(\Selector12~4_combout ),
	.datab(\Selector29~2_combout ),
	.datac(\ShiftLeft0~16_combout ),
	.datad(\Selector28~0_combout ),
	.cin(gnd),
	.combout(\Selector29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~3 .lut_mask = 16'h0800;
defparam \Selector29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N6
cycloneive_lcell_comb \ShiftRight0~74 (
// Equation(s):
// \ShiftRight0~74_combout  = (\portB~97_combout  & (\ShiftRight0~46_combout )) # (!\portB~97_combout  & ((\ShiftRight0~48_combout )))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftRight0~46_combout ),
	.datad(\ShiftRight0~48_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~74 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N12
cycloneive_lcell_comb \ShiftRight0~75 (
// Equation(s):
// \ShiftRight0~75_combout  = (\portB~100_combout  & (\ShiftRight0~45_combout  & (!\portB~97_combout ))) # (!\portB~100_combout  & (((\ShiftRight0~74_combout ))))

	.dataa(\ShiftRight0~45_combout ),
	.datab(portB30),
	.datac(portB31),
	.datad(\ShiftRight0~74_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~75 .lut_mask = 16'h2F20;
defparam \ShiftRight0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N26
cycloneive_lcell_comb \ShiftRight0~76 (
// Equation(s):
// \ShiftRight0~76_combout  = (\portB~97_combout  & ((\ShiftRight0~49_combout ))) # (!\portB~97_combout  & (\ShiftRight0~52_combout ))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftRight0~52_combout ),
	.datad(\ShiftRight0~49_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~76 .lut_mask = 16'hFC30;
defparam \ShiftRight0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N24
cycloneive_lcell_comb \ShiftRight0~55 (
// Equation(s):
// \ShiftRight0~55_combout  = (\portB~92_combout  & ((\portA~63_combout ))) # (!\portB~92_combout  & (\portA~65_combout ))

	.dataa(portA30),
	.datab(gnd),
	.datac(portA29),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~55 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N12
cycloneive_lcell_comb \ShiftRight0~77 (
// Equation(s):
// \ShiftRight0~77_combout  = (\portB~97_combout  & (\ShiftRight0~53_combout )) # (!\portB~97_combout  & ((\ShiftRight0~55_combout )))

	.dataa(\ShiftRight0~53_combout ),
	.datab(gnd),
	.datac(portB30),
	.datad(\ShiftRight0~55_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~77 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N6
cycloneive_lcell_comb \Selector21~0 (
// Equation(s):
// \Selector21~0_combout  = (\portB~100_combout  & (\ShiftRight0~76_combout )) # (!\portB~100_combout  & ((\ShiftRight0~77_combout )))

	.dataa(portB31),
	.datab(gnd),
	.datac(\ShiftRight0~76_combout ),
	.datad(\ShiftRight0~77_combout ),
	.cin(gnd),
	.combout(\Selector21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~0 .lut_mask = 16'hF5A0;
defparam \Selector21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N30
cycloneive_lcell_comb \ShiftRight0~78 (
// Equation(s):
// \ShiftRight0~78_combout  = (\portB~103_combout  & (\ShiftRight0~75_combout )) # (!\portB~103_combout  & ((\Selector21~0_combout )))

	.dataa(portB32),
	.datab(gnd),
	.datac(\ShiftRight0~75_combout ),
	.datad(\Selector21~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~78 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N30
cycloneive_lcell_comb \ShiftLeft0~20 (
// Equation(s):
// \ShiftLeft0~20_combout  = (!\portB~92_combout  & ((\portB~97_combout  & (\portA~69_combout )) # (!\portB~97_combout  & ((\portA~9_combout )))))

	.dataa(portB30),
	.datab(portA32),
	.datac(portA),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~20 .lut_mask = 16'h00D8;
defparam \ShiftLeft0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N24
cycloneive_lcell_comb \ShiftLeft0~21 (
// Equation(s):
// \ShiftLeft0~21_combout  = (\ShiftLeft0~20_combout ) # ((!\portB~97_combout  & (\portA~12_combout  & \portB~92_combout )))

	.dataa(portB30),
	.datab(portA1),
	.datac(\ShiftLeft0~20_combout ),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~21 .lut_mask = 16'hF4F0;
defparam \ShiftLeft0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N4
cycloneive_lcell_comb \Selector0~9 (
// Equation(s):
// \Selector0~9_combout  = (!ALUOp_EX[0] & (ALUOp_EX[2] & (!ALUOp_EX[3] & !ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~9 .lut_mask = 16'h0004;
defparam \Selector0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N28
cycloneive_lcell_comb \Selector29~4 (
// Equation(s):
// \Selector29~4_combout  = (\portA~9_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \portB~100_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(portA),
	.datad(portB31),
	.cin(gnd),
	.combout(\Selector29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~4 .lut_mask = 16'hE0A0;
defparam \Selector29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N10
cycloneive_lcell_comb \Selector29~5 (
// Equation(s):
// \Selector29~5_combout  = (\Selector29~4_combout ) # ((\Selector0~10_combout  & (\portB~100_combout  $ (\portA~9_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(portB31),
	.datac(portA),
	.datad(\Selector29~4_combout ),
	.cin(gnd),
	.combout(\Selector29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~5 .lut_mask = 16'hFF28;
defparam \Selector29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N22
cycloneive_lcell_comb \Selector29~6 (
// Equation(s):
// \Selector29~6_combout  = (\Selector0~13_combout  & (!\portA~9_combout  & !\portB~100_combout ))

	.dataa(gnd),
	.datab(\Selector0~13_combout ),
	.datac(portA),
	.datad(portB31),
	.cin(gnd),
	.combout(\Selector29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~6 .lut_mask = 16'h000C;
defparam \Selector29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N20
cycloneive_lcell_comb \Selector29~7 (
// Equation(s):
// \Selector29~7_combout  = (\Selector0~12_combout  & ((\Add0~4_combout ) # ((\Selector0~11_combout  & \Add1~4_combout )))) # (!\Selector0~12_combout  & (\Selector0~11_combout  & (\Add1~4_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Add1~4_combout ),
	.datad(\Add0~4_combout ),
	.cin(gnd),
	.combout(\Selector29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~7 .lut_mask = 16'hEAC0;
defparam \Selector29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N6
cycloneive_lcell_comb \Selector29~8 (
// Equation(s):
// \Selector29~8_combout  = (\Selector29~6_combout ) # ((\Selector29~7_combout ) # ((\Selector0~8_combout  & \portB~100_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(portB31),
	.datac(\Selector29~6_combout ),
	.datad(\Selector29~7_combout ),
	.cin(gnd),
	.combout(\Selector29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~8 .lut_mask = 16'hFFF8;
defparam \Selector29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N2
cycloneive_lcell_comb \Selector29~9 (
// Equation(s):
// \Selector29~9_combout  = (\Selector29~5_combout ) # ((\Selector29~8_combout ) # ((\ShiftLeft0~21_combout  & \Selector29~0_combout )))

	.dataa(\ShiftLeft0~21_combout ),
	.datab(\Selector29~5_combout ),
	.datac(\Selector29~0_combout ),
	.datad(\Selector29~8_combout ),
	.cin(gnd),
	.combout(\Selector29~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~9 .lut_mask = 16'hFFEC;
defparam \Selector29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N22
cycloneive_lcell_comb \Selector26~2 (
// Equation(s):
// \Selector26~2_combout  = (\portA~23_combout  & (((\Selector0~4_combout  & !\portB~87_combout )))) # (!\portA~23_combout  & ((\portB~87_combout  & ((\Selector0~4_combout ))) # (!\portB~87_combout  & (Selector0))))

	.dataa(Selector0),
	.datab(\Selector0~4_combout ),
	.datac(portA8),
	.datad(portB28),
	.cin(gnd),
	.combout(\Selector26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~2 .lut_mask = 16'h0CCA;
defparam \Selector26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N24
cycloneive_lcell_comb \Selector26~0 (
// Equation(s):
// \Selector26~0_combout  = (\Selector0~2_combout  & (((\portA~23_combout ) # (\portB~87_combout )))) # (!\Selector0~2_combout  & (\Selector0~3_combout  & (\portA~23_combout  & \portB~87_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(\Selector0~3_combout ),
	.datac(portA8),
	.datad(portB28),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~0 .lut_mask = 16'hEAA0;
defparam \Selector26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N8
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((\portA~14_combout  $ (\portB~107_combout  $ (\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((\portA~14_combout  & ((!\Add1~7 ) # (!\portB~107_combout ))) # (!\portA~14_combout  & (!\portB~107_combout  & !\Add1~7 )))

	.dataa(portA2),
	.datab(portB33),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h962B;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N10
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (\portA~23_combout  & ((\portB~87_combout  & (!\Add1~9 )) # (!\portB~87_combout  & (\Add1~9  & VCC)))) # (!\portA~23_combout  & ((\portB~87_combout  & ((\Add1~9 ) # (GND))) # (!\portB~87_combout  & (!\Add1~9 ))))
// \Add1~11  = CARRY((\portA~23_combout  & (\portB~87_combout  & !\Add1~9 )) # (!\portA~23_combout  & ((\portB~87_combout ) # (!\Add1~9 ))))

	.dataa(portA8),
	.datab(portB28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h694D;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N8
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = ((\portA~14_combout  $ (\portB~107_combout  $ (!\Add0~7 )))) # (GND)
// \Add0~9  = CARRY((\portA~14_combout  & ((\portB~107_combout ) # (!\Add0~7 ))) # (!\portA~14_combout  & (\portB~107_combout  & !\Add0~7 )))

	.dataa(portA2),
	.datab(portB33),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'h698E;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N10
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = (\portA~23_combout  & ((\portB~87_combout  & (\Add0~9  & VCC)) # (!\portB~87_combout  & (!\Add0~9 )))) # (!\portA~23_combout  & ((\portB~87_combout  & (!\Add0~9 )) # (!\portB~87_combout  & ((\Add0~9 ) # (GND)))))
// \Add0~11  = CARRY((\portA~23_combout  & (!\portB~87_combout  & !\Add0~9 )) # (!\portA~23_combout  & ((!\Add0~9 ) # (!\portB~87_combout ))))

	.dataa(portA8),
	.datab(portB28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h9617;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N12
cycloneive_lcell_comb \Selector26~1 (
// Equation(s):
// \Selector26~1_combout  = (\Add1~10_combout  & ((\Selector0~6_combout ) # ((\Selector0~7_combout  & \Add0~10_combout )))) # (!\Add1~10_combout  & (\Selector0~7_combout  & ((\Add0~10_combout ))))

	.dataa(\Add1~10_combout ),
	.datab(\Selector0~7_combout ),
	.datac(\Selector0~6_combout ),
	.datad(\Add0~10_combout ),
	.cin(gnd),
	.combout(\Selector26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~1 .lut_mask = 16'hECA0;
defparam \Selector26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N20
cycloneive_lcell_comb \Selector0~1 (
// Equation(s):
// \Selector0~1_combout  = (!ALUOp_EX[2] & (!ALUOp_EX[0] & (!ALUOp_EX[1] & !ALUOp_EX[3])))

	.dataa(ALUOp_EX_2),
	.datab(ALUOp_EX_0),
	.datac(ALUOp_EX_1),
	.datad(ALUOp_EX_3),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~1 .lut_mask = 16'h0001;
defparam \Selector0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N20
cycloneive_lcell_comb \Selector24~0 (
// Equation(s):
// \Selector24~0_combout  = (!\portB~103_combout  & (!\portB~107_combout  & (\Selector0~1_combout  & !\ShiftLeft0~16_combout )))

	.dataa(portB32),
	.datab(portB33),
	.datac(\Selector0~1_combout ),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~0 .lut_mask = 16'h0010;
defparam \Selector24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N12
cycloneive_lcell_comb \ShiftLeft0~22 (
// Equation(s):
// \ShiftLeft0~22_combout  = (\portB~92_combout  & ((\portA~14_combout ))) # (!\portB~92_combout  & (\portA~23_combout ))

	.dataa(portA8),
	.datab(portA2),
	.datac(portB29),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~22 .lut_mask = 16'hCACA;
defparam \ShiftLeft0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N6
cycloneive_lcell_comb \ShiftLeft0~23 (
// Equation(s):
// \ShiftLeft0~23_combout  = (\portB~97_combout  & (\ShiftLeft0~18_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~22_combout )))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftLeft0~18_combout ),
	.datad(\ShiftLeft0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~23 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N0
cycloneive_lcell_comb \ShiftLeft0~24 (
// Equation(s):
// \ShiftLeft0~24_combout  = (\portB~100_combout  & (!\portB~97_combout  & (\ShiftLeft0~13_combout ))) # (!\portB~100_combout  & (((\ShiftLeft0~23_combout ))))

	.dataa(portB30),
	.datab(portB31),
	.datac(\ShiftLeft0~13_combout ),
	.datad(\ShiftLeft0~23_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~24 .lut_mask = 16'h7340;
defparam \ShiftLeft0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N16
cycloneive_lcell_comb \Selector4~0 (
// Equation(s):
// \Selector4~0_combout  = (\portB~107_combout ) # ((!\portB~103_combout  & \portB~100_combout ))

	.dataa(gnd),
	.datab(portB32),
	.datac(portB33),
	.datad(portB31),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~0 .lut_mask = 16'hF3F0;
defparam \Selector4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N0
cycloneive_lcell_comb \ShiftRight0~80 (
// Equation(s):
// \ShiftRight0~80_combout  = (!\portB~103_combout  & ((\portB~100_combout  & (\ShiftRight0~21_combout )) # (!\portB~100_combout  & ((\ShiftRight0~25_combout )))))

	.dataa(portB31),
	.datab(portB32),
	.datac(\ShiftRight0~21_combout ),
	.datad(\ShiftRight0~25_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~80 .lut_mask = 16'h3120;
defparam \ShiftRight0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N22
cycloneive_lcell_comb \ShiftRight0~81 (
// Equation(s):
// \ShiftRight0~81_combout  = (\ShiftRight0~80_combout ) # ((\portB~103_combout  & (\ShiftRight0~18_combout  & !\portB~100_combout )))

	.dataa(portB32),
	.datab(\ShiftRight0~18_combout ),
	.datac(portB31),
	.datad(\ShiftRight0~80_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~81 .lut_mask = 16'hFF08;
defparam \ShiftRight0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N12
cycloneive_lcell_comb \ShiftRight0~11 (
// Equation(s):
// \ShiftRight0~11_combout  = (\portB~97_combout  & ((\ShiftRight0~9_combout ))) # (!\portB~97_combout  & (\ShiftRight0~10_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftRight0~10_combout ),
	.datad(\ShiftRight0~9_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~11 .lut_mask = 16'hFA50;
defparam \ShiftRight0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N10
cycloneive_lcell_comb \ShiftRight0~79 (
// Equation(s):
// \ShiftRight0~79_combout  = (\portB~100_combout  & (\ShiftRight0~28_combout )) # (!\portB~100_combout  & ((\ShiftRight0~11_combout )))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftRight0~28_combout ),
	.datad(\ShiftRight0~11_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~79 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N12
cycloneive_lcell_comb \Selector26~3 (
// Equation(s):
// \Selector26~3_combout  = (\Selector4~1_combout  & ((\Selector4~0_combout ) # ((\ShiftRight0~79_combout )))) # (!\Selector4~1_combout  & (!\Selector4~0_combout  & ((\ShiftRight0~7_combout ))))

	.dataa(\Selector4~1_combout ),
	.datab(\Selector4~0_combout ),
	.datac(\ShiftRight0~79_combout ),
	.datad(\ShiftRight0~7_combout ),
	.cin(gnd),
	.combout(\Selector26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~3 .lut_mask = 16'hB9A8;
defparam \Selector26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N2
cycloneive_lcell_comb \Selector26~4 (
// Equation(s):
// \Selector26~4_combout  = (\Selector4~0_combout  & ((\Selector26~3_combout  & ((\ShiftRight0~81_combout ))) # (!\Selector26~3_combout  & (\ShiftRight0~14_combout )))) # (!\Selector4~0_combout  & (((\Selector26~3_combout ))))

	.dataa(\ShiftRight0~14_combout ),
	.datab(\Selector4~0_combout ),
	.datac(\ShiftRight0~81_combout ),
	.datad(\Selector26~3_combout ),
	.cin(gnd),
	.combout(\Selector26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~4 .lut_mask = 16'hF388;
defparam \Selector26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N24
cycloneive_lcell_comb \Selector26~5 (
// Equation(s):
// \Selector26~5_combout  = (\Selector31~0_combout  & ((\Selector26~4_combout ) # ((\Selector24~0_combout  & \ShiftLeft0~24_combout )))) # (!\Selector31~0_combout  & (\Selector24~0_combout  & (\ShiftLeft0~24_combout )))

	.dataa(\Selector31~0_combout ),
	.datab(\Selector24~0_combout ),
	.datac(\ShiftLeft0~24_combout ),
	.datad(\Selector26~4_combout ),
	.cin(gnd),
	.combout(\Selector26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~5 .lut_mask = 16'hEAC0;
defparam \Selector26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N4
cycloneive_lcell_comb \ShiftLeft0~25 (
// Equation(s):
// \ShiftLeft0~25_combout  = (\portA~69_combout  & (!\portB~97_combout  & !\portB~92_combout ))

	.dataa(portA32),
	.datab(gnd),
	.datac(portB30),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~25 .lut_mask = 16'h000A;
defparam \ShiftLeft0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N2
cycloneive_lcell_comb \ShiftLeft0~27 (
// Equation(s):
// \ShiftLeft0~27_combout  = (\portB~92_combout  & (\portA~16_combout )) # (!\portB~92_combout  & ((\portA~14_combout )))

	.dataa(portA4),
	.datab(gnd),
	.datac(portA2),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~27 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N26
cycloneive_lcell_comb \ShiftLeft0~26 (
// Equation(s):
// \ShiftLeft0~26_combout  = (\portB~97_combout  & ((\portB~92_combout  & (\portA~12_combout )) # (!\portB~92_combout  & ((\portA~9_combout )))))

	.dataa(portB30),
	.datab(portA1),
	.datac(portA),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~26 .lut_mask = 16'h88A0;
defparam \ShiftLeft0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N8
cycloneive_lcell_comb \ShiftLeft0~28 (
// Equation(s):
// \ShiftLeft0~28_combout  = (\ShiftLeft0~26_combout ) # ((\ShiftLeft0~27_combout  & !\portB~97_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~27_combout ),
	.datac(portB30),
	.datad(\ShiftLeft0~26_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~28 .lut_mask = 16'hFF0C;
defparam \ShiftLeft0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N30
cycloneive_lcell_comb \ShiftLeft0~29 (
// Equation(s):
// \ShiftLeft0~29_combout  = (\portB~100_combout  & (\ShiftLeft0~25_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~28_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~25_combout ),
	.datac(\ShiftLeft0~28_combout ),
	.datad(portB31),
	.cin(gnd),
	.combout(\ShiftLeft0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~29 .lut_mask = 16'hCCF0;
defparam \ShiftLeft0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N26
cycloneive_lcell_comb \Selector4~1 (
// Equation(s):
// \Selector4~1_combout  = (\portB~107_combout ) # (\portB~103_combout )

	.dataa(gnd),
	.datab(portB33),
	.datac(portB32),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~1 .lut_mask = 16'hFCFC;
defparam \Selector4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N26
cycloneive_lcell_comb \ShiftRight0~56 (
// Equation(s):
// \ShiftRight0~56_combout  = (\portB~92_combout  & ((\portA~67_combout ))) # (!\portB~92_combout  & (\portA~25_combout ))

	.dataa(portA9),
	.datab(gnd),
	.datac(portA31),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~56 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N28
cycloneive_lcell_comb \ShiftRight0~57 (
// Equation(s):
// \ShiftRight0~57_combout  = (\portB~97_combout  & ((\ShiftRight0~55_combout ))) # (!\portB~97_combout  & (\ShiftRight0~56_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftRight0~56_combout ),
	.datad(\ShiftRight0~55_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~57 .lut_mask = 16'hFA50;
defparam \ShiftRight0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N30
cycloneive_lcell_comb \ShiftRight0~82 (
// Equation(s):
// \ShiftRight0~82_combout  = (\portB~100_combout  & (\ShiftRight0~57_combout )) # (!\portB~100_combout  & ((\ShiftRight0~39_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~57_combout ),
	.datac(portB31),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~82 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N4
cycloneive_lcell_comb \ShiftRight0~33 (
// Equation(s):
// \ShiftRight0~33_combout  = (\portB~92_combout  & (\portA~19_combout )) # (!\portB~92_combout  & ((\portA~21_combout )))

	.dataa(portA6),
	.datab(gnd),
	.datac(portA7),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftRight0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~33 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N26
cycloneive_lcell_comb \ShiftRight0~35 (
// Equation(s):
// \ShiftRight0~35_combout  = (\portB~97_combout  & (\ShiftRight0~33_combout )) # (!\portB~97_combout  & ((\ShiftRight0~34_combout )))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftRight0~33_combout ),
	.datad(\ShiftRight0~34_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~35 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N22
cycloneive_lcell_comb \Selector27~1 (
// Equation(s):
// \Selector27~1_combout  = (\Selector4~0_combout  & ((\ShiftRight0~42_combout ) # ((\Selector4~1_combout )))) # (!\Selector4~0_combout  & (((!\Selector4~1_combout  & \ShiftRight0~35_combout ))))

	.dataa(\Selector4~0_combout ),
	.datab(\ShiftRight0~42_combout ),
	.datac(\Selector4~1_combout ),
	.datad(\ShiftRight0~35_combout ),
	.cin(gnd),
	.combout(\Selector27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~1 .lut_mask = 16'hADA8;
defparam \Selector27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N16
cycloneive_lcell_comb \ShiftRight0~83 (
// Equation(s):
// \ShiftRight0~83_combout  = (!\portB~103_combout  & ((\portB~100_combout  & (\ShiftRight0~50_combout )) # (!\portB~100_combout  & ((\ShiftRight0~54_combout )))))

	.dataa(portB32),
	.datab(portB31),
	.datac(\ShiftRight0~50_combout ),
	.datad(\ShiftRight0~54_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~83 .lut_mask = 16'h5140;
defparam \ShiftRight0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N18
cycloneive_lcell_comb \ShiftRight0~84 (
// Equation(s):
// \ShiftRight0~84_combout  = (\ShiftRight0~83_combout ) # ((\portB~103_combout  & (\ShiftRight0~47_combout  & !\portB~100_combout )))

	.dataa(portB32),
	.datab(\ShiftRight0~47_combout ),
	.datac(portB31),
	.datad(\ShiftRight0~83_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~84 .lut_mask = 16'hFF08;
defparam \ShiftRight0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N16
cycloneive_lcell_comb \Selector27~2 (
// Equation(s):
// \Selector27~2_combout  = (\Selector4~1_combout  & ((\Selector27~1_combout  & ((\ShiftRight0~84_combout ))) # (!\Selector27~1_combout  & (\ShiftRight0~82_combout )))) # (!\Selector4~1_combout  & (((\Selector27~1_combout ))))

	.dataa(\Selector4~1_combout ),
	.datab(\ShiftRight0~82_combout ),
	.datac(\Selector27~1_combout ),
	.datad(\ShiftRight0~84_combout ),
	.cin(gnd),
	.combout(\Selector27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~2 .lut_mask = 16'hF858;
defparam \Selector27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N2
cycloneive_lcell_comb \Selector27~4 (
// Equation(s):
// \Selector27~4_combout  = (\portA~14_combout  & ((\Selector0~3_combout ))) # (!\portA~14_combout  & (Selector0))

	.dataa(Selector0),
	.datab(portA2),
	.datac(gnd),
	.datad(\Selector0~3_combout ),
	.cin(gnd),
	.combout(\Selector27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~4 .lut_mask = 16'hEE22;
defparam \Selector27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N0
cycloneive_lcell_comb \Selector27~5 (
// Equation(s):
// \Selector27~5_combout  = (\portB~107_combout  & ((\Selector0~2_combout ) # (!\portA~14_combout ))) # (!\portB~107_combout  & ((\portA~14_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(gnd),
	.datac(portB33),
	.datad(portA2),
	.cin(gnd),
	.combout(\Selector27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~5 .lut_mask = 16'hAFF0;
defparam \Selector27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N14
cycloneive_lcell_comb \ShiftRight0~85 (
// Equation(s):
// \ShiftRight0~85_combout  = (\portB~100_combout  & (\ShiftRight0~68_combout )) # (!\portB~100_combout  & ((\ShiftRight0~60_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~68_combout ),
	.datac(\ShiftRight0~60_combout ),
	.datad(portB31),
	.cin(gnd),
	.combout(\ShiftRight0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~85 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N18
cycloneive_lcell_comb \Selector24~6 (
// Equation(s):
// \Selector24~6_combout  = (\Selector4~1_combout  & (((\Selector4~0_combout )))) # (!\Selector4~1_combout  & ((\Selector4~0_combout  & (\ShiftRight0~61_combout )) # (!\Selector4~0_combout  & ((\ShiftRight0~59_combout )))))

	.dataa(\ShiftRight0~61_combout ),
	.datab(\Selector4~1_combout ),
	.datac(\ShiftRight0~59_combout ),
	.datad(\Selector4~0_combout ),
	.cin(gnd),
	.combout(\Selector24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~6 .lut_mask = 16'hEE30;
defparam \Selector24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N16
cycloneive_lcell_comb \Selector24~7 (
// Equation(s):
// \Selector24~7_combout  = (\Selector4~1_combout  & ((\Selector24~6_combout  & ((ShiftRight0))) # (!\Selector24~6_combout  & (\ShiftRight0~85_combout )))) # (!\Selector4~1_combout  & (((\Selector24~6_combout ))))

	.dataa(\Selector4~1_combout ),
	.datab(\ShiftRight0~85_combout ),
	.datac(ShiftRight0),
	.datad(\Selector24~6_combout ),
	.cin(gnd),
	.combout(\Selector24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~7 .lut_mask = 16'hF588;
defparam \Selector24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N28
cycloneive_lcell_comb \Selector24~1 (
// Equation(s):
// \Selector24~1_combout  = (\portA~19_combout  & ((\Selector0~2_combout ) # ((\Selector0~3_combout  & \portB~82_combout )))) # (!\portA~19_combout  & (((\portB~82_combout  & \Selector0~2_combout ))))

	.dataa(portA6),
	.datab(\Selector0~3_combout ),
	.datac(portB26),
	.datad(\Selector0~2_combout ),
	.cin(gnd),
	.combout(\Selector24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~1 .lut_mask = 16'hFA80;
defparam \Selector24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N22
cycloneive_lcell_comb \Selector24~3 (
// Equation(s):
// \Selector24~3_combout  = (\portB~82_combout  & (\Selector0~4_combout  & ((!\portA~19_combout )))) # (!\portB~82_combout  & ((\portA~19_combout  & (\Selector0~4_combout )) # (!\portA~19_combout  & ((Selector0)))))

	.dataa(portB26),
	.datab(\Selector0~4_combout ),
	.datac(Selector0),
	.datad(portA6),
	.cin(gnd),
	.combout(\Selector24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~3 .lut_mask = 16'h44D8;
defparam \Selector24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N14
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (\portA~19_combout  & ((\portB~82_combout  & (!\Add1~13 )) # (!\portB~82_combout  & (\Add1~13  & VCC)))) # (!\portA~19_combout  & ((\portB~82_combout  & ((\Add1~13 ) # (GND))) # (!\portB~82_combout  & (!\Add1~13 ))))
// \Add1~15  = CARRY((\portA~19_combout  & (\portB~82_combout  & !\Add1~13 )) # (!\portA~19_combout  & ((\portB~82_combout ) # (!\Add1~13 ))))

	.dataa(portA6),
	.datab(portB26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h694D;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N12
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = ((\portA~21_combout  $ (\portB~84_combout  $ (!\Add0~11 )))) # (GND)
// \Add0~13  = CARRY((\portA~21_combout  & ((\portB~84_combout ) # (!\Add0~11 ))) # (!\portA~21_combout  & (\portB~84_combout  & !\Add0~11 )))

	.dataa(portA7),
	.datab(portB27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'h698E;
defparam \Add0~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N14
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = (\portB~82_combout  & ((\portA~19_combout  & (\Add0~13  & VCC)) # (!\portA~19_combout  & (!\Add0~13 )))) # (!\portB~82_combout  & ((\portA~19_combout  & (!\Add0~13 )) # (!\portA~19_combout  & ((\Add0~13 ) # (GND)))))
// \Add0~15  = CARRY((\portB~82_combout  & (!\portA~19_combout  & !\Add0~13 )) # (!\portB~82_combout  & ((!\Add0~13 ) # (!\portA~19_combout ))))

	.dataa(portB26),
	.datab(portA6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h9617;
defparam \Add0~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N10
cycloneive_lcell_comb \Selector24~2 (
// Equation(s):
// \Selector24~2_combout  = (\Selector0~7_combout  & ((\Add0~14_combout ) # ((\Selector0~6_combout  & \Add1~14_combout )))) # (!\Selector0~7_combout  & (\Selector0~6_combout  & (\Add1~14_combout )))

	.dataa(\Selector0~7_combout ),
	.datab(\Selector0~6_combout ),
	.datac(\Add1~14_combout ),
	.datad(\Add0~14_combout ),
	.cin(gnd),
	.combout(\Selector24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~2 .lut_mask = 16'hEAC0;
defparam \Selector24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N8
cycloneive_lcell_comb \Selector24~4 (
// Equation(s):
// \Selector24~4_combout  = (\Selector24~1_combout ) # ((\Selector24~3_combout ) # (\Selector24~2_combout ))

	.dataa(gnd),
	.datab(\Selector24~1_combout ),
	.datac(\Selector24~3_combout ),
	.datad(\Selector24~2_combout ),
	.cin(gnd),
	.combout(\Selector24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~4 .lut_mask = 16'hFFFC;
defparam \Selector24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N30
cycloneive_lcell_comb \ShiftLeft0~30 (
// Equation(s):
// \ShiftLeft0~30_combout  = (\portB~92_combout  & ((\portA~21_combout ))) # (!\portB~92_combout  & (\portA~19_combout ))

	.dataa(portA6),
	.datab(gnd),
	.datac(portB29),
	.datad(portA7),
	.cin(gnd),
	.combout(\ShiftLeft0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~30 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N16
cycloneive_lcell_comb \ShiftLeft0~31 (
// Equation(s):
// \ShiftLeft0~31_combout  = (\portB~97_combout  & ((\ShiftLeft0~22_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~30_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftLeft0~30_combout ),
	.datad(\ShiftLeft0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~31 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N18
cycloneive_lcell_comb \ShiftLeft0~32 (
// Equation(s):
// \ShiftLeft0~32_combout  = (\portB~100_combout  & (\ShiftLeft0~19_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~31_combout )))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftLeft0~19_combout ),
	.datad(\ShiftLeft0~31_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~32 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N10
cycloneive_lcell_comb \Selector4~2 (
// Equation(s):
// \Selector4~2_combout  = (\ShiftLeft0~12_combout ) # ((\portB~103_combout ) # ((\portB~107_combout ) # (\ShiftLeft0~6_combout )))

	.dataa(\ShiftLeft0~12_combout ),
	.datab(portB32),
	.datac(portB33),
	.datad(\ShiftLeft0~6_combout ),
	.cin(gnd),
	.combout(\Selector4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~2 .lut_mask = 16'hFFFE;
defparam \Selector4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N2
cycloneive_lcell_comb \Selector24~5 (
// Equation(s):
// \Selector24~5_combout  = (\Selector0~1_combout  & (\ShiftLeft0~32_combout  & !\Selector4~2_combout ))

	.dataa(\Selector0~1_combout ),
	.datab(\ShiftLeft0~32_combout ),
	.datac(\Selector4~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~5 .lut_mask = 16'h0808;
defparam \Selector24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N12
cycloneive_lcell_comb \Selector25~2 (
// Equation(s):
// \Selector25~2_combout  = (\portA~21_combout  & (((\Selector0~4_combout  & !\portB~84_combout )))) # (!\portA~21_combout  & ((\portB~84_combout  & ((\Selector0~4_combout ))) # (!\portB~84_combout  & (Selector0))))

	.dataa(Selector0),
	.datab(\Selector0~4_combout ),
	.datac(portA7),
	.datad(portB27),
	.cin(gnd),
	.combout(\Selector25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~2 .lut_mask = 16'h0CCA;
defparam \Selector25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N30
cycloneive_lcell_comb \Selector25~0 (
// Equation(s):
// \Selector25~0_combout  = (\Selector0~2_combout  & (((\portA~21_combout ) # (\portB~84_combout )))) # (!\Selector0~2_combout  & (\Selector0~3_combout  & (\portA~21_combout  & \portB~84_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(\Selector0~3_combout ),
	.datac(portA7),
	.datad(portB27),
	.cin(gnd),
	.combout(\Selector25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~0 .lut_mask = 16'hEAA0;
defparam \Selector25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N16
cycloneive_lcell_comb \Selector25~1 (
// Equation(s):
// \Selector25~1_combout  = (\Add1~12_combout  & ((\Selector0~6_combout ) # ((\Selector0~7_combout  & \Add0~12_combout )))) # (!\Add1~12_combout  & (\Selector0~7_combout  & ((\Add0~12_combout ))))

	.dataa(\Add1~12_combout ),
	.datab(\Selector0~7_combout ),
	.datac(\Selector0~6_combout ),
	.datad(\Add0~12_combout ),
	.cin(gnd),
	.combout(\Selector25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~1 .lut_mask = 16'hECA0;
defparam \Selector25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N26
cycloneive_lcell_comb \Selector25~3 (
// Equation(s):
// \Selector25~3_combout  = (\Selector25~2_combout ) # ((\Selector25~0_combout ) # (\Selector25~1_combout ))

	.dataa(gnd),
	.datab(\Selector25~2_combout ),
	.datac(\Selector25~0_combout ),
	.datad(\Selector25~1_combout ),
	.cin(gnd),
	.combout(\Selector25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~3 .lut_mask = 16'hFFFC;
defparam \Selector25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N2
cycloneive_lcell_comb \ShiftRight0~89 (
// Equation(s):
// \ShiftRight0~89_combout  = (\ShiftRight0~45_combout  & (!\portB~97_combout  & (!\portB~100_combout  & \portB~103_combout )))

	.dataa(\ShiftRight0~45_combout ),
	.datab(portB30),
	.datac(portB31),
	.datad(portB32),
	.cin(gnd),
	.combout(\ShiftRight0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~89 .lut_mask = 16'h0200;
defparam \ShiftRight0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N28
cycloneive_lcell_comb \Selector4~3 (
// Equation(s):
// \Selector4~3_combout  = (!\portB~103_combout  & \portB~100_combout )

	.dataa(portB32),
	.datab(gnd),
	.datac(portB31),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~3 .lut_mask = 16'h5050;
defparam \Selector4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N2
cycloneive_lcell_comb \ShiftRight0~88 (
// Equation(s):
// \ShiftRight0~88_combout  = (\Selector4~3_combout  & ((\portB~97_combout  & (\ShiftRight0~46_combout )) # (!\portB~97_combout  & ((\ShiftRight0~48_combout )))))

	.dataa(portB30),
	.datab(\ShiftRight0~46_combout ),
	.datac(\ShiftRight0~48_combout ),
	.datad(\Selector4~3_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~88 .lut_mask = 16'hD800;
defparam \ShiftRight0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N30
cycloneive_lcell_comb \ShiftRight0~90 (
// Equation(s):
// \ShiftRight0~90_combout  = (\ShiftRight0~89_combout ) # ((\ShiftRight0~88_combout ) # ((\ShiftRight0~76_combout  & \ShiftLeft0~17_combout )))

	.dataa(\ShiftRight0~76_combout ),
	.datab(\ShiftRight0~89_combout ),
	.datac(\ShiftLeft0~17_combout ),
	.datad(\ShiftRight0~88_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~90 .lut_mask = 16'hFFEC;
defparam \ShiftRight0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N4
cycloneive_lcell_comb \ShiftRight0~87 (
// Equation(s):
// \ShiftRight0~87_combout  = (\portB~100_combout  & (\ShiftRight0~77_combout )) # (!\portB~100_combout  & ((\ShiftRight0~71_combout )))

	.dataa(\ShiftRight0~77_combout ),
	.datab(gnd),
	.datac(portB31),
	.datad(\ShiftRight0~71_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~87 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N18
cycloneive_lcell_comb \Selector25~5 (
// Equation(s):
// \Selector25~5_combout  = (\Selector4~1_combout  & (((\ShiftRight0~87_combout ) # (\Selector4~0_combout )))) # (!\Selector4~1_combout  & (\ShiftRight0~70_combout  & ((!\Selector4~0_combout ))))

	.dataa(\ShiftRight0~70_combout ),
	.datab(\ShiftRight0~87_combout ),
	.datac(\Selector4~1_combout ),
	.datad(\Selector4~0_combout ),
	.cin(gnd),
	.combout(\Selector25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~5 .lut_mask = 16'hF0CA;
defparam \Selector25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N20
cycloneive_lcell_comb \Selector25~6 (
// Equation(s):
// \Selector25~6_combout  = (\Selector4~0_combout  & ((\Selector25~5_combout  & (\ShiftRight0~90_combout )) # (!\Selector25~5_combout  & ((\ShiftRight0~72_combout ))))) # (!\Selector4~0_combout  & (((\Selector25~5_combout ))))

	.dataa(\ShiftRight0~90_combout ),
	.datab(\ShiftRight0~72_combout ),
	.datac(\Selector4~0_combout ),
	.datad(\Selector25~5_combout ),
	.cin(gnd),
	.combout(\Selector25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~6 .lut_mask = 16'hAFC0;
defparam \Selector25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N0
cycloneive_lcell_comb \ShiftLeft0~35 (
// Equation(s):
// \ShiftLeft0~35_combout  = (\portB~100_combout  & ((\ShiftLeft0~21_combout ))) # (!\portB~100_combout  & (\ShiftLeft0~34_combout ))

	.dataa(\ShiftLeft0~34_combout ),
	.datab(\ShiftLeft0~21_combout ),
	.datac(gnd),
	.datad(portB31),
	.cin(gnd),
	.combout(\ShiftLeft0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~35 .lut_mask = 16'hCCAA;
defparam \ShiftLeft0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N28
cycloneive_lcell_comb \Selector25~4 (
// Equation(s):
// \Selector25~4_combout  = (\Selector0~1_combout  & (\ShiftLeft0~35_combout  & !\Selector4~2_combout ))

	.dataa(gnd),
	.datab(\Selector0~1_combout ),
	.datac(\ShiftLeft0~35_combout ),
	.datad(\Selector4~2_combout ),
	.cin(gnd),
	.combout(\Selector25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~4 .lut_mask = 16'h00C0;
defparam \Selector25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N0
cycloneive_lcell_comb \Selector0~12 (
// Equation(s):
// \Selector0~12_combout  = (!ALUOp_EX[0] & (!ALUOp_EX[2] & (!ALUOp_EX[3] & ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~12 .lut_mask = 16'h0100;
defparam \Selector0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N16
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = ((\portA~17_combout  $ (\portB~76_combout  $ (!\Add0~15 )))) # (GND)
// \Add0~17  = CARRY((\portA~17_combout  & ((\portB~76_combout ) # (!\Add0~15 ))) # (!\portA~17_combout  & (\portB~76_combout  & !\Add0~15 )))

	.dataa(portA5),
	.datab(portB23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'h698E;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N18
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = (\portB~73_combout  & ((\portA~37_combout  & (\Add0~17  & VCC)) # (!\portA~37_combout  & (!\Add0~17 )))) # (!\portB~73_combout  & ((\portA~37_combout  & (!\Add0~17 )) # (!\portA~37_combout  & ((\Add0~17 ) # (GND)))))
// \Add0~19  = CARRY((\portB~73_combout  & (!\portA~37_combout  & !\Add0~17 )) # (!\portB~73_combout  & ((!\Add0~17 ) # (!\portA~37_combout ))))

	.dataa(portB21),
	.datab(portA16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h9617;
defparam \Add0~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N26
cycloneive_lcell_comb \Selector22~7 (
// Equation(s):
// \Selector22~7_combout  = (\Selector0~12_combout  & \Add0~18_combout )

	.dataa(\Selector0~12_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Add0~18_combout ),
	.cin(gnd),
	.combout(\Selector22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~7 .lut_mask = 16'hAA00;
defparam \Selector22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N16
cycloneive_lcell_comb \ShiftLeft0~38 (
// Equation(s):
// \ShiftLeft0~38_combout  = (\portB~92_combout  & (\portA~17_combout )) # (!\portB~92_combout  & ((\portA~37_combout )))

	.dataa(portA5),
	.datab(gnd),
	.datac(portA16),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~38 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N20
cycloneive_lcell_comb \ShiftLeft0~39 (
// Equation(s):
// \ShiftLeft0~39_combout  = (\portB~97_combout  & (\ShiftLeft0~30_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~38_combout )))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftLeft0~30_combout ),
	.datad(\ShiftLeft0~38_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~39 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N4
cycloneive_lcell_comb \ShiftLeft0~36 (
// Equation(s):
// \ShiftLeft0~36_combout  = (\Selector4~3_combout  & ((\portB~97_combout  & (\ShiftLeft0~18_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~22_combout )))))

	.dataa(portB30),
	.datab(\ShiftLeft0~18_combout ),
	.datac(\ShiftLeft0~22_combout ),
	.datad(\Selector4~3_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~36 .lut_mask = 16'hD800;
defparam \ShiftLeft0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N22
cycloneive_lcell_comb \ShiftLeft0~40 (
// Equation(s):
// \ShiftLeft0~40_combout  = (\ShiftLeft0~37_combout ) # ((\ShiftLeft0~36_combout ) # ((\ShiftLeft0~39_combout  & \ShiftLeft0~17_combout )))

	.dataa(\ShiftLeft0~37_combout ),
	.datab(\ShiftLeft0~39_combout ),
	.datac(\ShiftLeft0~36_combout ),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~40 .lut_mask = 16'hFEFA;
defparam \ShiftLeft0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N14
cycloneive_lcell_comb \Selector22~5 (
// Equation(s):
// \Selector22~5_combout  = (\Selector0~14_combout  & (!\portB~107_combout  & (!\ShiftLeft0~16_combout  & \ShiftLeft0~40_combout )))

	.dataa(\Selector0~14_combout ),
	.datab(portB33),
	.datac(\ShiftLeft0~16_combout ),
	.datad(\ShiftLeft0~40_combout ),
	.cin(gnd),
	.combout(\Selector22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~5 .lut_mask = 16'h0200;
defparam \Selector22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N18
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (\portB~73_combout  & ((\portA~37_combout  & (!\Add1~17 )) # (!\portA~37_combout  & ((\Add1~17 ) # (GND))))) # (!\portB~73_combout  & ((\portA~37_combout  & (\Add1~17  & VCC)) # (!\portA~37_combout  & (!\Add1~17 ))))
// \Add1~19  = CARRY((\portB~73_combout  & ((!\Add1~17 ) # (!\portA~37_combout ))) # (!\portB~73_combout  & (!\portA~37_combout  & !\Add1~17 )))

	.dataa(portB21),
	.datab(portA16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h692B;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N24
cycloneive_lcell_comb \Selector22~6 (
// Equation(s):
// \Selector22~6_combout  = (\Selector22~5_combout ) # ((\Selector0~11_combout  & \Add1~18_combout ))

	.dataa(\Selector0~11_combout ),
	.datab(\Selector22~5_combout ),
	.datac(gnd),
	.datad(\Add1~18_combout ),
	.cin(gnd),
	.combout(\Selector22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~6 .lut_mask = 16'hEECC;
defparam \Selector22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N30
cycloneive_lcell_comb \Selector22~3 (
// Equation(s):
// \Selector22~3_combout  = (\Selector0~8_combout  & (((\portA~37_combout ) # (\portB~73_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\portA~37_combout  & \portB~73_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(portA16),
	.datad(portB21),
	.cin(gnd),
	.combout(\Selector22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~3 .lut_mask = 16'hEAA0;
defparam \Selector22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N20
cycloneive_lcell_comb \Selector22~2 (
// Equation(s):
// \Selector22~2_combout  = (\portA~37_combout  & (\Selector0~10_combout  & ((!\portB~73_combout )))) # (!\portA~37_combout  & ((\portB~73_combout  & (\Selector0~10_combout )) # (!\portB~73_combout  & ((\Selector0~13_combout )))))

	.dataa(portA16),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~13_combout ),
	.datad(portB21),
	.cin(gnd),
	.combout(\Selector22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~2 .lut_mask = 16'h44D8;
defparam \Selector22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N18
cycloneive_lcell_comb \Selector16~1 (
// Equation(s):
// \Selector16~1_combout  = (ALUOp_EX[0] & ((\ShiftLeft0~16_combout ) # ((!\portB~103_combout  & !\portB~107_combout ))))

	.dataa(ALUOp_EX_0),
	.datab(portB32),
	.datac(portB33),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~1 .lut_mask = 16'hAA02;
defparam \Selector16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N6
cycloneive_lcell_comb \Selector16~2 (
// Equation(s):
// \Selector16~2_combout  = (\Selector12~5_combout  & \Selector16~1_combout )

	.dataa(gnd),
	.datab(\Selector12~5_combout ),
	.datac(gnd),
	.datad(\Selector16~1_combout ),
	.cin(gnd),
	.combout(\Selector16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~2 .lut_mask = 16'hCC00;
defparam \Selector16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N4
cycloneive_lcell_comb \Selector22~4 (
// Equation(s):
// \Selector22~4_combout  = (\Selector22~3_combout ) # ((\Selector22~2_combout ) # ((\Selector16~2_combout  & \ShiftRight0~15_combout )))

	.dataa(\Selector22~3_combout ),
	.datab(\Selector22~2_combout ),
	.datac(\Selector16~2_combout ),
	.datad(\ShiftRight0~15_combout ),
	.cin(gnd),
	.combout(\Selector22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~4 .lut_mask = 16'hFEEE;
defparam \Selector22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N6
cycloneive_lcell_comb \Selector20~1 (
// Equation(s):
// \Selector20~1_combout  = (!\portB~103_combout  & (ALUOp_EX[0] & (\portB~107_combout  & \Selector12~5_combout )))

	.dataa(portB32),
	.datab(ALUOp_EX_0),
	.datac(portB33),
	.datad(\Selector12~5_combout ),
	.cin(gnd),
	.combout(\Selector20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~1 .lut_mask = 16'h4000;
defparam \Selector20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N0
cycloneive_lcell_comb \Selector12~6 (
// Equation(s):
// \Selector12~6_combout  = (\portB~103_combout  & (ALUOp_EX[0] & (!\portB~107_combout  & \Selector12~5_combout )))

	.dataa(portB32),
	.datab(ALUOp_EX_0),
	.datac(portB33),
	.datad(\Selector12~5_combout ),
	.cin(gnd),
	.combout(\Selector12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~6 .lut_mask = 16'h0800;
defparam \Selector12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N8
cycloneive_lcell_comb \Selector22~1 (
// Equation(s):
// \Selector22~1_combout  = (\ShiftRight0~22_combout  & ((\Selector20~1_combout ) # ((\Selector12~6_combout  & \Selector22~0_combout )))) # (!\ShiftRight0~22_combout  & (((\Selector12~6_combout  & \Selector22~0_combout ))))

	.dataa(\ShiftRight0~22_combout ),
	.datab(\Selector20~1_combout ),
	.datac(\Selector12~6_combout ),
	.datad(\Selector22~0_combout ),
	.cin(gnd),
	.combout(\Selector22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~1 .lut_mask = 16'hF888;
defparam \Selector22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N18
cycloneive_lcell_comb \Selector0~14 (
// Equation(s):
// \Selector0~14_combout  = (!ALUOp_EX[0] & (!ALUOp_EX[2] & (!ALUOp_EX[3] & !ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~14 .lut_mask = 16'h0001;
defparam \Selector0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N6
cycloneive_lcell_comb \ShiftLeft0~41 (
// Equation(s):
// \ShiftLeft0~41_combout  = (\portB~103_combout  & (\ShiftLeft0~25_combout  & ((!\portB~100_combout )))) # (!\portB~103_combout  & (((\ShiftLeft0~28_combout  & \portB~100_combout ))))

	.dataa(\ShiftLeft0~25_combout ),
	.datab(portB32),
	.datac(\ShiftLeft0~28_combout ),
	.datad(portB31),
	.cin(gnd),
	.combout(\ShiftLeft0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~41 .lut_mask = 16'h3088;
defparam \ShiftLeft0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N10
cycloneive_lcell_comb \ShiftLeft0~42 (
// Equation(s):
// \ShiftLeft0~42_combout  = (\portB~92_combout  & ((\portA~19_combout ))) # (!\portB~92_combout  & (\portA~17_combout ))

	.dataa(portA5),
	.datab(gnd),
	.datac(portA6),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~42 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N12
cycloneive_lcell_comb \ShiftLeft0~33 (
// Equation(s):
// \ShiftLeft0~33_combout  = (\portB~92_combout  & ((\portA~23_combout ))) # (!\portB~92_combout  & (\portA~21_combout ))

	.dataa(gnd),
	.datab(portA7),
	.datac(portA8),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~33 .lut_mask = 16'hF0CC;
defparam \ShiftLeft0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N18
cycloneive_lcell_comb \ShiftLeft0~43 (
// Equation(s):
// \ShiftLeft0~43_combout  = (\portB~97_combout  & ((\ShiftLeft0~33_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~42_combout ))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftLeft0~42_combout ),
	.datad(\ShiftLeft0~33_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~43 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N26
cycloneive_lcell_comb \Selector23~1 (
// Equation(s):
// \Selector23~1_combout  = (Selector16 & ((\ShiftLeft0~41_combout ) # ((\ShiftLeft0~17_combout  & \ShiftLeft0~43_combout ))))

	.dataa(\ShiftLeft0~17_combout ),
	.datab(\ShiftLeft0~41_combout ),
	.datac(\ShiftLeft0~43_combout ),
	.datad(Selector16),
	.cin(gnd),
	.combout(\Selector23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~1 .lut_mask = 16'hEC00;
defparam \Selector23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N4
cycloneive_lcell_comb \Selector23~3 (
// Equation(s):
// \Selector23~3_combout  = (\portA~17_combout ) # ((\portB~76_combout ) # (\Selector0~13_combout ))

	.dataa(portA5),
	.datab(gnd),
	.datac(portB23),
	.datad(\Selector0~13_combout ),
	.cin(gnd),
	.combout(\Selector23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~3 .lut_mask = 16'hFFFA;
defparam \Selector23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N12
cycloneive_lcell_comb \Selector23~2 (
// Equation(s):
// \Selector23~2_combout  = (\portA~17_combout  & ((\portB~76_combout  & ((\Selector0~9_combout ))) # (!\portB~76_combout  & (\Selector0~10_combout )))) # (!\portA~17_combout  & ((\Selector0~10_combout ) # ((!\portB~76_combout ))))

	.dataa(portA5),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~9_combout ),
	.datad(portB23),
	.cin(gnd),
	.combout(\Selector23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~2 .lut_mask = 16'hE4DD;
defparam \Selector23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N8
cycloneive_lcell_comb \Selector23~4 (
// Equation(s):
// \Selector23~4_combout  = (\Selector23~3_combout  & ((\Selector0~8_combout ) # (\Selector23~2_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(gnd),
	.datac(\Selector23~3_combout ),
	.datad(\Selector23~2_combout ),
	.cin(gnd),
	.combout(\Selector23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~4 .lut_mask = 16'hF0A0;
defparam \Selector23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N30
cycloneive_lcell_comb \Selector23~5 (
// Equation(s):
// \Selector23~5_combout  = (\Selector23~4_combout ) # ((\Selector23~0_combout  & \Selector12~6_combout ))

	.dataa(gnd),
	.datab(\Selector23~0_combout ),
	.datac(\Selector23~4_combout ),
	.datad(\Selector12~6_combout ),
	.cin(gnd),
	.combout(\Selector23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~5 .lut_mask = 16'hFCF0;
defparam \Selector23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N20
cycloneive_lcell_comb \Selector23~6 (
// Equation(s):
// \Selector23~6_combout  = (\Add1~16_combout  & ((\Selector0~11_combout ) # ((\Selector16~2_combout  & \ShiftRight0~43_combout )))) # (!\Add1~16_combout  & (((\Selector16~2_combout  & \ShiftRight0~43_combout ))))

	.dataa(\Add1~16_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Selector16~2_combout ),
	.datad(\ShiftRight0~43_combout ),
	.cin(gnd),
	.combout(\Selector23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~6 .lut_mask = 16'hF888;
defparam \Selector23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N18
cycloneive_lcell_comb \Selector23~7 (
// Equation(s):
// \Selector23~7_combout  = (\Selector23~5_combout ) # ((\Selector23~6_combout ) # ((\Add0~16_combout  & \Selector0~12_combout )))

	.dataa(\Add0~16_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Selector23~5_combout ),
	.datad(\Selector23~6_combout ),
	.cin(gnd),
	.combout(\Selector23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~7 .lut_mask = 16'hFFF8;
defparam \Selector23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N20
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = ((\portA~36_combout  $ (\portB~109_combout  $ (!\Add0~19 )))) # (GND)
// \Add0~21  = CARRY((\portA~36_combout  & ((\portB~109_combout ) # (!\Add0~19 ))) # (!\portA~36_combout  & (\portB~109_combout  & !\Add0~19 )))

	.dataa(portA15),
	.datab(portB35),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'h698E;
defparam \Add0~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N22
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = (\portA~35_combout  & ((\portB~108_combout  & (\Add0~21  & VCC)) # (!\portB~108_combout  & (!\Add0~21 )))) # (!\portA~35_combout  & ((\portB~108_combout  & (!\Add0~21 )) # (!\portB~108_combout  & ((\Add0~21 ) # (GND)))))
// \Add0~23  = CARRY((\portA~35_combout  & (!\portB~108_combout  & !\Add0~21 )) # (!\portA~35_combout  & ((!\Add0~21 ) # (!\portB~108_combout ))))

	.dataa(portA14),
	.datab(portB34),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h9617;
defparam \Add0~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N20
cycloneive_lcell_comb \Selector20~2 (
// Equation(s):
// \Selector20~2_combout  = (\portA~35_combout  & (\Selector0~10_combout  & ((!\portB~108_combout )))) # (!\portA~35_combout  & ((\portB~108_combout  & (\Selector0~10_combout )) # (!\portB~108_combout  & ((\Selector0~13_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~13_combout ),
	.datac(portA14),
	.datad(portB34),
	.cin(gnd),
	.combout(\Selector20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~2 .lut_mask = 16'h0AAC;
defparam \Selector20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N4
cycloneive_lcell_comb \Selector20~3 (
// Equation(s):
// \Selector20~3_combout  = (\ShiftLeft0~47_combout  & ((Selector16) # ((\Selector20~0_combout  & \Selector12~6_combout )))) # (!\ShiftLeft0~47_combout  & (((\Selector20~0_combout  & \Selector12~6_combout ))))

	.dataa(\ShiftLeft0~47_combout ),
	.datab(Selector16),
	.datac(\Selector20~0_combout ),
	.datad(\Selector12~6_combout ),
	.cin(gnd),
	.combout(\Selector20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~3 .lut_mask = 16'hF888;
defparam \Selector20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N20
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((\portB~109_combout  $ (\portA~36_combout  $ (\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((\portB~109_combout  & (\portA~36_combout  & !\Add1~19 )) # (!\portB~109_combout  & ((\portA~36_combout ) # (!\Add1~19 ))))

	.dataa(portB35),
	.datab(portA15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h964D;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N22
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (\portA~35_combout  & ((\portB~108_combout  & (!\Add1~21 )) # (!\portB~108_combout  & (\Add1~21  & VCC)))) # (!\portA~35_combout  & ((\portB~108_combout  & ((\Add1~21 ) # (GND))) # (!\portB~108_combout  & (!\Add1~21 ))))
// \Add1~23  = CARRY((\portA~35_combout  & (\portB~108_combout  & !\Add1~21 )) # (!\portA~35_combout  & ((\portB~108_combout ) # (!\Add1~21 ))))

	.dataa(portA14),
	.datab(portB34),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h694D;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N14
cycloneive_lcell_comb \Selector20~4 (
// Equation(s):
// \Selector20~4_combout  = (\Selector20~2_combout ) # ((\Selector20~3_combout ) # ((\Selector0~11_combout  & \Add1~22_combout )))

	.dataa(\Selector20~2_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Selector20~3_combout ),
	.datad(\Add1~22_combout ),
	.cin(gnd),
	.combout(\Selector20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~4 .lut_mask = 16'hFEFA;
defparam \Selector20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N26
cycloneive_lcell_comb \Selector20~5 (
// Equation(s):
// \Selector20~5_combout  = (\portA~35_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \portB~108_combout )))) # (!\portA~35_combout  & (\Selector0~8_combout  & ((\portB~108_combout ))))

	.dataa(portA14),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~9_combout ),
	.datad(portB34),
	.cin(gnd),
	.combout(\Selector20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~5 .lut_mask = 16'hEC88;
defparam \Selector20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N8
cycloneive_lcell_comb \Selector20~6 (
// Equation(s):
// \Selector20~6_combout  = (\ShiftRight0~66_combout  & ((\Selector20~1_combout ) # ((\ShiftRight0~62_combout  & \Selector16~2_combout )))) # (!\ShiftRight0~66_combout  & (\ShiftRight0~62_combout  & ((\Selector16~2_combout ))))

	.dataa(\ShiftRight0~66_combout ),
	.datab(\ShiftRight0~62_combout ),
	.datac(\Selector20~1_combout ),
	.datad(\Selector16~2_combout ),
	.cin(gnd),
	.combout(\Selector20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~6 .lut_mask = 16'hECA0;
defparam \Selector20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N28
cycloneive_lcell_comb \Selector20~7 (
// Equation(s):
// \Selector20~7_combout  = (\Selector20~5_combout ) # (\Selector20~6_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Selector20~5_combout ),
	.datad(\Selector20~6_combout ),
	.cin(gnd),
	.combout(\Selector20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~7 .lut_mask = 16'hFFF0;
defparam \Selector20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N24
cycloneive_lcell_comb \Selector21~4 (
// Equation(s):
// \Selector21~4_combout  = (\portA~36_combout  & (\Selector0~10_combout  & (!\portB~109_combout ))) # (!\portA~36_combout  & ((\portB~109_combout  & (\Selector0~10_combout )) # (!\portB~109_combout  & ((\Selector0~13_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(portA15),
	.datac(portB35),
	.datad(\Selector0~13_combout ),
	.cin(gnd),
	.combout(\Selector21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~4 .lut_mask = 16'h2B28;
defparam \Selector21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N6
cycloneive_lcell_comb \ShiftLeft0~34 (
// Equation(s):
// \ShiftLeft0~34_combout  = (\portB~97_combout  & (\ShiftLeft0~27_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~33_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~27_combout ),
	.datac(portB30),
	.datad(\ShiftLeft0~33_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~34 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N4
cycloneive_lcell_comb \ShiftLeft0~48 (
// Equation(s):
// \ShiftLeft0~48_combout  = (\portB~92_combout  & (\portA~37_combout )) # (!\portB~92_combout  & ((\portA~36_combout )))

	.dataa(portA16),
	.datab(gnd),
	.datac(portA15),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~48 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N22
cycloneive_lcell_comb \ShiftLeft0~49 (
// Equation(s):
// \ShiftLeft0~49_combout  = (\portB~97_combout  & ((\ShiftLeft0~42_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~48_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftLeft0~48_combout ),
	.datad(\ShiftLeft0~42_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~49 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N12
cycloneive_lcell_comb \ShiftLeft0~50 (
// Equation(s):
// \ShiftLeft0~50_combout  = (!\portB~103_combout  & ((\portB~100_combout  & (\ShiftLeft0~34_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~49_combout )))))

	.dataa(portB32),
	.datab(portB31),
	.datac(\ShiftLeft0~34_combout ),
	.datad(\ShiftLeft0~49_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~50 .lut_mask = 16'h5140;
defparam \ShiftLeft0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N18
cycloneive_lcell_comb \ShiftLeft0~51 (
// Equation(s):
// \ShiftLeft0~51_combout  = (\ShiftLeft0~50_combout ) # ((\portB~103_combout  & (!\portB~100_combout  & \ShiftLeft0~21_combout )))

	.dataa(portB32),
	.datab(portB31),
	.datac(\ShiftLeft0~21_combout ),
	.datad(\ShiftLeft0~50_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~51 .lut_mask = 16'hFF20;
defparam \ShiftLeft0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N0
cycloneive_lcell_comb \Selector21~5 (
// Equation(s):
// \Selector21~5_combout  = (\Selector21~3_combout ) # ((\Selector21~4_combout ) # ((Selector16 & \ShiftLeft0~51_combout )))

	.dataa(\Selector21~3_combout ),
	.datab(Selector16),
	.datac(\Selector21~4_combout ),
	.datad(\ShiftLeft0~51_combout ),
	.cin(gnd),
	.combout(\Selector21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~5 .lut_mask = 16'hFEFA;
defparam \Selector21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N2
cycloneive_lcell_comb \Selector21~2 (
// Equation(s):
// \Selector21~2_combout  = (\Selector12~5_combout  & (\ShiftRight0~73_combout  & \Selector16~1_combout ))

	.dataa(gnd),
	.datab(\Selector12~5_combout ),
	.datac(\ShiftRight0~73_combout ),
	.datad(\Selector16~1_combout ),
	.cin(gnd),
	.combout(\Selector21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~2 .lut_mask = 16'hC000;
defparam \Selector21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N14
cycloneive_lcell_comb \Selector21~6 (
// Equation(s):
// \Selector21~6_combout  = (\Selector21~5_combout ) # ((\Selector21~2_combout ) # ((\Selector0~11_combout  & \Add1~20_combout )))

	.dataa(\Selector0~11_combout ),
	.datab(\Selector21~5_combout ),
	.datac(\Add1~20_combout ),
	.datad(\Selector21~2_combout ),
	.cin(gnd),
	.combout(\Selector21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~6 .lut_mask = 16'hFFEC;
defparam \Selector21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N2
cycloneive_lcell_comb \Selector21~1 (
// Equation(s):
// \Selector21~1_combout  = (\Selector21~0_combout  & ((\Selector12~6_combout ) # ((\ShiftRight0~75_combout  & \Selector20~1_combout )))) # (!\Selector21~0_combout  & (((\ShiftRight0~75_combout  & \Selector20~1_combout ))))

	.dataa(\Selector21~0_combout ),
	.datab(\Selector12~6_combout ),
	.datac(\ShiftRight0~75_combout ),
	.datad(\Selector20~1_combout ),
	.cin(gnd),
	.combout(\Selector21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~1 .lut_mask = 16'hF888;
defparam \Selector21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N30
cycloneive_lcell_comb \Selector18~0 (
// Equation(s):
// \Selector18~0_combout  = (!\portB~103_combout  & (\Selector16~0_combout  & (!\portB~100_combout  & \ShiftRight0~18_combout )))

	.dataa(portB32),
	.datab(\Selector16~0_combout ),
	.datac(portB31),
	.datad(\ShiftRight0~18_combout ),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~0 .lut_mask = 16'h0400;
defparam \Selector18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N30
cycloneive_lcell_comb \Selector18~2 (
// Equation(s):
// \Selector18~2_combout  = (\portA~31_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \portB~68_combout )))) # (!\portA~31_combout  & (((\portB~68_combout  & \Selector0~8_combout ))))

	.dataa(\Selector0~9_combout ),
	.datab(portA12),
	.datac(portB18),
	.datad(\Selector0~8_combout ),
	.cin(gnd),
	.combout(\Selector18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~2 .lut_mask = 16'hFC80;
defparam \Selector18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N4
cycloneive_lcell_comb \Selector18~3 (
// Equation(s):
// \Selector18~3_combout  = (\portB~68_combout  & (\Selector0~10_combout  & ((!\portA~31_combout )))) # (!\portB~68_combout  & ((\portA~31_combout  & (\Selector0~10_combout )) # (!\portA~31_combout  & ((\Selector0~13_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~13_combout ),
	.datac(portB18),
	.datad(portA12),
	.cin(gnd),
	.combout(\Selector18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~3 .lut_mask = 16'h0AAC;
defparam \Selector18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N24
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((\portA~33_combout  $ (\portB~70_combout  $ (\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((\portA~33_combout  & ((!\Add1~23 ) # (!\portB~70_combout ))) # (!\portA~33_combout  & (!\portB~70_combout  & !\Add1~23 )))

	.dataa(portA13),
	.datab(portB19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h962B;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N26
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (\portA~31_combout  & ((\portB~68_combout  & (!\Add1~25 )) # (!\portB~68_combout  & (\Add1~25  & VCC)))) # (!\portA~31_combout  & ((\portB~68_combout  & ((\Add1~25 ) # (GND))) # (!\portB~68_combout  & (!\Add1~25 ))))
// \Add1~27  = CARRY((\portA~31_combout  & (\portB~68_combout  & !\Add1~25 )) # (!\portA~31_combout  & ((\portB~68_combout ) # (!\Add1~25 ))))

	.dataa(portA12),
	.datab(portB18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h694D;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N14
cycloneive_lcell_comb \Selector18~4 (
// Equation(s):
// \Selector18~4_combout  = (\Selector18~2_combout ) # ((\Selector18~3_combout ) # ((\Selector0~11_combout  & \Add1~26_combout )))

	.dataa(\Selector18~2_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Selector18~3_combout ),
	.datad(\Add1~26_combout ),
	.cin(gnd),
	.combout(\Selector18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~4 .lut_mask = 16'hFEFA;
defparam \Selector18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N20
cycloneive_lcell_comb \ShiftLeft0~52 (
// Equation(s):
// \ShiftLeft0~52_combout  = (\portB~92_combout  & (\portA~33_combout )) # (!\portB~92_combout  & ((\portA~31_combout )))

	.dataa(portA13),
	.datab(gnd),
	.datac(portA12),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~52 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N12
cycloneive_lcell_comb \ShiftLeft0~44 (
// Equation(s):
// \ShiftLeft0~44_combout  = (\portB~92_combout  & (\portA~36_combout )) # (!\portB~92_combout  & ((\portA~35_combout )))

	.dataa(gnd),
	.datab(portA15),
	.datac(portB29),
	.datad(portA14),
	.cin(gnd),
	.combout(\ShiftLeft0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~44 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N18
cycloneive_lcell_comb \ShiftLeft0~53 (
// Equation(s):
// \ShiftLeft0~53_combout  = (\portB~97_combout  & ((\ShiftLeft0~44_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~52_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~52_combout ),
	.datac(portB30),
	.datad(\ShiftLeft0~44_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~53 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N8
cycloneive_lcell_comb \Selector10~0 (
// Equation(s):
// \Selector10~0_combout  = (\portB~100_combout  & ((\ShiftLeft0~39_combout ))) # (!\portB~100_combout  & (\ShiftLeft0~53_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~53_combout ),
	.datac(portB31),
	.datad(\ShiftLeft0~39_combout ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~0 .lut_mask = 16'hFC0C;
defparam \Selector10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N26
cycloneive_lcell_comb \ShiftLeft0~54 (
// Equation(s):
// \ShiftLeft0~54_combout  = (\portB~103_combout  & ((\ShiftLeft0~24_combout ))) # (!\portB~103_combout  & (\Selector10~0_combout ))

	.dataa(portB32),
	.datab(gnd),
	.datac(\Selector10~0_combout ),
	.datad(\ShiftLeft0~24_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~54 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N28
cycloneive_lcell_comb \Selector18~1 (
// Equation(s):
// \Selector18~1_combout  = (\Selector16~2_combout  & ((\ShiftRight0~79_combout ) # ((Selector16 & \ShiftLeft0~54_combout )))) # (!\Selector16~2_combout  & (Selector16 & ((\ShiftLeft0~54_combout ))))

	.dataa(\Selector16~2_combout ),
	.datab(Selector16),
	.datac(\ShiftRight0~79_combout ),
	.datad(\ShiftLeft0~54_combout ),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~1 .lut_mask = 16'hECA0;
defparam \Selector18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N24
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = ((\portB~70_combout  $ (\portA~33_combout  $ (!\Add0~23 )))) # (GND)
// \Add0~25  = CARRY((\portB~70_combout  & ((\portA~33_combout ) # (!\Add0~23 ))) # (!\portB~70_combout  & (\portA~33_combout  & !\Add0~23 )))

	.dataa(portB19),
	.datab(portA13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'h698E;
defparam \Add0~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N26
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = (\portA~31_combout  & ((\portB~68_combout  & (\Add0~25  & VCC)) # (!\portB~68_combout  & (!\Add0~25 )))) # (!\portA~31_combout  & ((\portB~68_combout  & (!\Add0~25 )) # (!\portB~68_combout  & ((\Add0~25 ) # (GND)))))
// \Add0~27  = CARRY((\portA~31_combout  & (!\portB~68_combout  & !\Add0~25 )) # (!\portA~31_combout  & ((!\Add0~25 ) # (!\portB~68_combout ))))

	.dataa(portA12),
	.datab(portB18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h9617;
defparam \Add0~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N4
cycloneive_lcell_comb \Selector18~5 (
// Equation(s):
// \Selector18~5_combout  = (\Selector12~6_combout  & ((\portB~100_combout  & (\ShiftRight0~21_combout )) # (!\portB~100_combout  & ((\ShiftRight0~25_combout )))))

	.dataa(\ShiftRight0~21_combout ),
	.datab(portB31),
	.datac(\ShiftRight0~25_combout ),
	.datad(\Selector12~6_combout ),
	.cin(gnd),
	.combout(\Selector18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~5 .lut_mask = 16'hB800;
defparam \Selector18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N12
cycloneive_lcell_comb \Selector18~6 (
// Equation(s):
// \Selector18~6_combout  = (\Selector18~5_combout ) # ((\Selector0~12_combout  & \Add0~26_combout ))

	.dataa(\Selector0~12_combout ),
	.datab(gnd),
	.datac(\Add0~26_combout ),
	.datad(\Selector18~5_combout ),
	.cin(gnd),
	.combout(\Selector18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~6 .lut_mask = 16'hFFA0;
defparam \Selector18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N0
cycloneive_lcell_comb \Selector19~3 (
// Equation(s):
// \Selector19~3_combout  = (\portB~70_combout  & (\Selector0~10_combout  & ((!\portA~33_combout )))) # (!\portB~70_combout  & ((\portA~33_combout  & (\Selector0~10_combout )) # (!\portA~33_combout  & ((\Selector0~13_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~13_combout ),
	.datac(portB19),
	.datad(portA13),
	.cin(gnd),
	.combout(\Selector19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~3 .lut_mask = 16'h0AAC;
defparam \Selector19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N8
cycloneive_lcell_comb \Selector19~4 (
// Equation(s):
// \Selector19~4_combout  = (\Selector19~3_combout ) # ((\ShiftLeft0~17_combout  & (\ShiftRight0~47_combout  & \Selector16~0_combout )))

	.dataa(\ShiftLeft0~17_combout ),
	.datab(\Selector19~3_combout ),
	.datac(\ShiftRight0~47_combout ),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~4 .lut_mask = 16'hECCC;
defparam \Selector19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N26
cycloneive_lcell_comb \Selector19~5 (
// Equation(s):
// \Selector19~5_combout  = (\Selector19~4_combout ) # ((\Selector0~11_combout  & \Add1~24_combout ))

	.dataa(\Selector0~11_combout ),
	.datab(gnd),
	.datac(\Selector19~4_combout ),
	.datad(\Add1~24_combout ),
	.cin(gnd),
	.combout(\Selector19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~5 .lut_mask = 16'hFAF0;
defparam \Selector19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N10
cycloneive_lcell_comb \Selector19~0 (
// Equation(s):
// \Selector19~0_combout  = (\portA~33_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \portB~70_combout )))) # (!\portA~33_combout  & (((\portB~70_combout  & \Selector0~8_combout ))))

	.dataa(portA13),
	.datab(\Selector0~9_combout ),
	.datac(portB19),
	.datad(\Selector0~8_combout ),
	.cin(gnd),
	.combout(\Selector19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~0 .lut_mask = 16'hFA80;
defparam \Selector19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N10
cycloneive_lcell_comb \Selector19~1 (
// Equation(s):
// \Selector19~1_combout  = (\Selector12~6_combout  & ((\portB~100_combout  & ((\ShiftRight0~50_combout ))) # (!\portB~100_combout  & (\ShiftRight0~54_combout ))))

	.dataa(portB31),
	.datab(\ShiftRight0~54_combout ),
	.datac(\ShiftRight0~50_combout ),
	.datad(\Selector12~6_combout ),
	.cin(gnd),
	.combout(\Selector19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~1 .lut_mask = 16'hE400;
defparam \Selector19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N10
cycloneive_lcell_comb \Selector19~2 (
// Equation(s):
// \Selector19~2_combout  = (\Selector19~0_combout ) # ((\Selector19~1_combout ) # ((\Selector16~2_combout  & \ShiftRight0~82_combout )))

	.dataa(\Selector16~2_combout ),
	.datab(\ShiftRight0~82_combout ),
	.datac(\Selector19~0_combout ),
	.datad(\Selector19~1_combout ),
	.cin(gnd),
	.combout(\Selector19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~2 .lut_mask = 16'hFFF8;
defparam \Selector19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N16
cycloneive_lcell_comb \ShiftLeft0~55 (
// Equation(s):
// \ShiftLeft0~55_combout  = (\portB~92_combout  & (\portA~35_combout )) # (!\portB~92_combout  & ((\portA~33_combout )))

	.dataa(portA14),
	.datab(gnd),
	.datac(portA13),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~55 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N22
cycloneive_lcell_comb \ShiftLeft0~56 (
// Equation(s):
// \ShiftLeft0~56_combout  = (\portB~97_combout  & (\ShiftLeft0~48_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~55_combout )))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftLeft0~48_combout ),
	.datad(\ShiftLeft0~55_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~56 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N20
cycloneive_lcell_comb \Selector11~0 (
// Equation(s):
// \Selector11~0_combout  = (\portB~100_combout  & ((\ShiftLeft0~43_combout ))) # (!\portB~100_combout  & (\ShiftLeft0~56_combout ))

	.dataa(portB31),
	.datab(gnd),
	.datac(\ShiftLeft0~56_combout ),
	.datad(\ShiftLeft0~43_combout ),
	.cin(gnd),
	.combout(\Selector11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~0 .lut_mask = 16'hFA50;
defparam \Selector11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N28
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = ((\portB~66_combout  $ (\portA~29_combout  $ (!\Add0~27 )))) # (GND)
// \Add0~29  = CARRY((\portB~66_combout  & ((\portA~29_combout ) # (!\Add0~27 ))) # (!\portB~66_combout  & (\portA~29_combout  & !\Add0~27 )))

	.dataa(portB17),
	.datab(portA11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'h698E;
defparam \Add0~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N30
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = (\portB~64_combout  & ((\portA~27_combout  & (\Add0~29  & VCC)) # (!\portA~27_combout  & (!\Add0~29 )))) # (!\portB~64_combout  & ((\portA~27_combout  & (!\Add0~29 )) # (!\portA~27_combout  & ((\Add0~29 ) # (GND)))))
// \Add0~31  = CARRY((\portB~64_combout  & (!\portA~27_combout  & !\Add0~29 )) # (!\portB~64_combout  & ((!\Add0~29 ) # (!\portA~27_combout ))))

	.dataa(portB16),
	.datab(portA10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h9617;
defparam \Add0~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N12
cycloneive_lcell_comb \Selector16~4 (
// Equation(s):
// \Selector16~4_combout  = (\portA~27_combout  & (\Selector0~10_combout  & (!\portB~64_combout ))) # (!\portA~27_combout  & ((\portB~64_combout  & (\Selector0~10_combout )) # (!\portB~64_combout  & ((\Selector0~13_combout )))))

	.dataa(portA10),
	.datab(\Selector0~10_combout ),
	.datac(portB16),
	.datad(\Selector0~13_combout ),
	.cin(gnd),
	.combout(\Selector16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~4 .lut_mask = 16'h4D48;
defparam \Selector16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N12
cycloneive_lcell_comb \Selector16~5 (
// Equation(s):
// \Selector16~5_combout  = (\Selector12~6_combout  & ((\portB~100_combout  & (\ShiftRight0~65_combout )) # (!\portB~100_combout  & ((\ShiftRight0~67_combout )))))

	.dataa(\ShiftRight0~65_combout ),
	.datab(portB31),
	.datac(\ShiftRight0~67_combout ),
	.datad(\Selector12~6_combout ),
	.cin(gnd),
	.combout(\Selector16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~5 .lut_mask = 16'hB800;
defparam \Selector16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N8
cycloneive_lcell_comb \Selector16~6 (
// Equation(s):
// \Selector16~6_combout  = (\portA~39_combout  & (!\ShiftLeft0~15_combout  & \Selector16~0_combout ))

	.dataa(gnd),
	.datab(portA17),
	.datac(\ShiftLeft0~15_combout ),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~6 .lut_mask = 16'h0C00;
defparam \Selector16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N26
cycloneive_lcell_comb \ShiftLeft0~58 (
// Equation(s):
// \ShiftLeft0~58_combout  = (\portB~92_combout  & ((\portA~29_combout ))) # (!\portB~92_combout  & (\portA~27_combout ))

	.dataa(portA10),
	.datab(portA11),
	.datac(gnd),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~58 .lut_mask = 16'hCCAA;
defparam \ShiftLeft0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N4
cycloneive_lcell_comb \ShiftLeft0~59 (
// Equation(s):
// \ShiftLeft0~59_combout  = (\portB~97_combout  & ((\ShiftLeft0~52_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~58_combout ))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftLeft0~58_combout ),
	.datad(\ShiftLeft0~52_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~59 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N6
cycloneive_lcell_comb \ShiftLeft0~45 (
// Equation(s):
// \ShiftLeft0~45_combout  = (\portB~97_combout  & (\ShiftLeft0~38_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~44_combout )))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftLeft0~38_combout ),
	.datad(\ShiftLeft0~44_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~45 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N2
cycloneive_lcell_comb \Selector8~0 (
// Equation(s):
// \Selector8~0_combout  = (\portB~100_combout  & ((\ShiftLeft0~45_combout ))) # (!\portB~100_combout  & (\ShiftLeft0~59_combout ))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftLeft0~59_combout ),
	.datad(\ShiftLeft0~45_combout ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~0 .lut_mask = 16'hFC30;
defparam \Selector8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N22
cycloneive_lcell_comb \ShiftLeft0~60 (
// Equation(s):
// \ShiftLeft0~60_combout  = (\portB~103_combout  & (\ShiftLeft0~32_combout )) # (!\portB~103_combout  & ((\Selector8~0_combout )))

	.dataa(gnd),
	.datab(portB32),
	.datac(\ShiftLeft0~32_combout ),
	.datad(\Selector8~0_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~60 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N16
cycloneive_lcell_comb \Selector16~7 (
// Equation(s):
// \Selector16~7_combout  = (Selector16 & ((\ShiftLeft0~60_combout ) # ((\ShiftRight0~85_combout  & \Selector16~2_combout )))) # (!Selector16 & (\ShiftRight0~85_combout  & ((\Selector16~2_combout ))))

	.dataa(Selector16),
	.datab(\ShiftRight0~85_combout ),
	.datac(\ShiftLeft0~60_combout ),
	.datad(\Selector16~2_combout ),
	.cin(gnd),
	.combout(\Selector16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~7 .lut_mask = 16'hECA0;
defparam \Selector16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N26
cycloneive_lcell_comb \Selector16~8 (
// Equation(s):
// \Selector16~8_combout  = (\Selector16~4_combout ) # ((\Selector16~5_combout ) # ((\Selector16~6_combout ) # (\Selector16~7_combout )))

	.dataa(\Selector16~4_combout ),
	.datab(\Selector16~5_combout ),
	.datac(\Selector16~6_combout ),
	.datad(\Selector16~7_combout ),
	.cin(gnd),
	.combout(\Selector16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~8 .lut_mask = 16'hFFFE;
defparam \Selector16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N14
cycloneive_lcell_comb \Selector16~9 (
// Equation(s):
// \Selector16~9_combout  = (\Selector0~8_combout  & (((\portB~64_combout ) # (\portA~27_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\portB~64_combout  & \portA~27_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector0~8_combout ),
	.datac(portB16),
	.datad(portA10),
	.cin(gnd),
	.combout(\Selector16~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~9 .lut_mask = 16'hECC0;
defparam \Selector16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N28
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((\portA~29_combout  $ (\portB~66_combout  $ (\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((\portA~29_combout  & ((!\Add1~27 ) # (!\portB~66_combout ))) # (!\portA~29_combout  & (!\portB~66_combout  & !\Add1~27 )))

	.dataa(portA11),
	.datab(portB17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h962B;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N30
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (\portA~27_combout  & ((\portB~64_combout  & (!\Add1~29 )) # (!\portB~64_combout  & (\Add1~29  & VCC)))) # (!\portA~27_combout  & ((\portB~64_combout  & ((\Add1~29 ) # (GND))) # (!\portB~64_combout  & (!\Add1~29 ))))
// \Add1~31  = CARRY((\portA~27_combout  & (\portB~64_combout  & !\Add1~29 )) # (!\portA~27_combout  & ((\portB~64_combout ) # (!\Add1~29 ))))

	.dataa(portA10),
	.datab(portB16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h694D;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N28
cycloneive_lcell_comb \Selector16~10 (
// Equation(s):
// \Selector16~10_combout  = (\Selector16~9_combout ) # ((\Selector0~11_combout  & \Add1~30_combout ))

	.dataa(gnd),
	.datab(\Selector0~11_combout ),
	.datac(\Selector16~9_combout ),
	.datad(\Add1~30_combout ),
	.cin(gnd),
	.combout(\Selector16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~10 .lut_mask = 16'hFCF0;
defparam \Selector16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N22
cycloneive_lcell_comb \Selector17~9 (
// Equation(s):
// \Selector17~9_combout  = (!\portB~97_combout  & (!\portB~100_combout  & (\ShiftRight0~45_combout  & \Selector20~1_combout )))

	.dataa(portB30),
	.datab(portB31),
	.datac(\ShiftRight0~45_combout ),
	.datad(\Selector20~1_combout ),
	.cin(gnd),
	.combout(\Selector17~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~9 .lut_mask = 16'h1000;
defparam \Selector17~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N4
cycloneive_lcell_comb \ShiftLeft0~61 (
// Equation(s):
// \ShiftLeft0~61_combout  = (\portB~92_combout  & (\portA~31_combout )) # (!\portB~92_combout  & ((\portA~29_combout )))

	.dataa(gnd),
	.datab(portA12),
	.datac(portA11),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~61 .lut_mask = 16'hCCF0;
defparam \ShiftLeft0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N28
cycloneive_lcell_comb \ShiftLeft0~62 (
// Equation(s):
// \ShiftLeft0~62_combout  = (\portB~97_combout  & ((\ShiftLeft0~55_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~61_combout ))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftLeft0~61_combout ),
	.datad(\ShiftLeft0~55_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~62 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N22
cycloneive_lcell_comb \Selector9~0 (
// Equation(s):
// \Selector9~0_combout  = (\portB~100_combout  & (\ShiftLeft0~49_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~62_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~49_combout ),
	.datac(portB31),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~0 .lut_mask = 16'hCFC0;
defparam \Selector9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N26
cycloneive_lcell_comb \ShiftLeft0~63 (
// Equation(s):
// \ShiftLeft0~63_combout  = (\portB~103_combout  & (\ShiftLeft0~35_combout )) # (!\portB~103_combout  & ((\Selector9~0_combout )))

	.dataa(gnd),
	.datab(portB32),
	.datac(\ShiftLeft0~35_combout ),
	.datad(\Selector9~0_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~63 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N8
cycloneive_lcell_comb \Selector17~2 (
// Equation(s):
// \Selector17~2_combout  = (Selector16 & ((\ShiftLeft0~63_combout ) # ((\ShiftRight0~87_combout  & \Selector16~2_combout )))) # (!Selector16 & (\ShiftRight0~87_combout  & ((\Selector16~2_combout ))))

	.dataa(Selector16),
	.datab(\ShiftRight0~87_combout ),
	.datac(\ShiftLeft0~63_combout ),
	.datad(\Selector16~2_combout ),
	.cin(gnd),
	.combout(\Selector17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~2 .lut_mask = 16'hECA0;
defparam \Selector17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N16
cycloneive_lcell_comb \Selector17~4 (
// Equation(s):
// \Selector17~4_combout  = (\portB~66_combout  & (\Selector0~10_combout  & ((!\portA~29_combout )))) # (!\portB~66_combout  & ((\portA~29_combout  & (\Selector0~10_combout )) # (!\portA~29_combout  & ((\Selector0~13_combout )))))

	.dataa(portB17),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~13_combout ),
	.datad(portA11),
	.cin(gnd),
	.combout(\Selector17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~4 .lut_mask = 16'h44D8;
defparam \Selector17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N18
cycloneive_lcell_comb \Selector17~3 (
// Equation(s):
// \Selector17~3_combout  = (\portB~66_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \portA~29_combout )))) # (!\portB~66_combout  & (\Selector0~8_combout  & ((\portA~29_combout ))))

	.dataa(portB17),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~9_combout ),
	.datad(portA11),
	.cin(gnd),
	.combout(\Selector17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~3 .lut_mask = 16'hEC88;
defparam \Selector17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N6
cycloneive_lcell_comb \Selector17~5 (
// Equation(s):
// \Selector17~5_combout  = (\Selector17~4_combout ) # ((\Selector17~3_combout ) # ((\Selector0~11_combout  & \Add1~28_combout )))

	.dataa(\Selector0~11_combout ),
	.datab(\Selector17~4_combout ),
	.datac(\Add1~28_combout ),
	.datad(\Selector17~3_combout ),
	.cin(gnd),
	.combout(\Selector17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~5 .lut_mask = 16'hFFEC;
defparam \Selector17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N18
cycloneive_lcell_comb \Selector17~6 (
// Equation(s):
// \Selector17~6_combout  = (\Selector12~6_combout  & ((\portB~100_combout  & (\ShiftRight0~74_combout )) # (!\portB~100_combout  & ((\ShiftRight0~76_combout )))))

	.dataa(\ShiftRight0~74_combout ),
	.datab(portB31),
	.datac(\Selector12~6_combout ),
	.datad(\ShiftRight0~76_combout ),
	.cin(gnd),
	.combout(\Selector17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~6 .lut_mask = 16'hB080;
defparam \Selector17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N24
cycloneive_lcell_comb \Selector17~7 (
// Equation(s):
// \Selector17~7_combout  = (\Selector17~6_combout ) # ((\Selector0~12_combout  & \Add0~28_combout ))

	.dataa(\Selector0~12_combout ),
	.datab(\Add0~28_combout ),
	.datac(gnd),
	.datad(\Selector17~6_combout ),
	.cin(gnd),
	.combout(\Selector17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~7 .lut_mask = 16'hFF88;
defparam \Selector17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N8
cycloneive_lcell_comb \Selector0~15 (
// Equation(s):
// \Selector0~15_combout  = (ALUOp_EX[0] & (!ALUOp_EX[2] & (!ALUOp_EX[3] & !ALUOp_EX[1])))

	.dataa(ALUOp_EX_0),
	.datab(ALUOp_EX_2),
	.datac(ALUOp_EX_3),
	.datad(ALUOp_EX_1),
	.cin(gnd),
	.combout(\Selector0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~15 .lut_mask = 16'h0002;
defparam \Selector0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N0
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_combout  = ((\portB~62_combout  $ (\portA~25_combout  $ (!\Add0~31 )))) # (GND)
// \Add0~33  = CARRY((\portB~62_combout  & ((\portA~25_combout ) # (!\Add0~31 ))) # (!\portB~62_combout  & (\portA~25_combout  & !\Add0~31 )))

	.dataa(portB15),
	.datab(portA9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'h698E;
defparam \Add0~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N2
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = (\portA~67_combout  & ((\portB~59_combout  & (\Add0~33  & VCC)) # (!\portB~59_combout  & (!\Add0~33 )))) # (!\portA~67_combout  & ((\portB~59_combout  & (!\Add0~33 )) # (!\portB~59_combout  & ((\Add0~33 ) # (GND)))))
// \Add0~35  = CARRY((\portA~67_combout  & (!\portB~59_combout  & !\Add0~33 )) # (!\portA~67_combout  & ((!\Add0~33 ) # (!\portB~59_combout ))))

	.dataa(portA31),
	.datab(portB14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout(\Add0~35 ));
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h9617;
defparam \Add0~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N10
cycloneive_lcell_comb \Selector14~1 (
// Equation(s):
// \Selector14~1_combout  = (\portB~59_combout  & (\Selector0~10_combout  & ((!\portA~67_combout )))) # (!\portB~59_combout  & ((\portA~67_combout  & (\Selector0~10_combout )) # (!\portA~67_combout  & ((\Selector0~13_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~13_combout ),
	.datac(portB14),
	.datad(portA31),
	.cin(gnd),
	.combout(\Selector14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~1 .lut_mask = 16'h0AAC;
defparam \Selector14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N18
cycloneive_lcell_comb \Selector14~0 (
// Equation(s):
// \Selector14~0_combout  = (\portA~67_combout  & ((\Selector0~8_combout ) # ((\portB~59_combout  & \Selector0~9_combout )))) # (!\portA~67_combout  & (\Selector0~8_combout  & (\portB~59_combout )))

	.dataa(portA31),
	.datab(\Selector0~8_combout ),
	.datac(portB14),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~0 .lut_mask = 16'hE8C8;
defparam \Selector14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N24
cycloneive_lcell_comb \Selector12~7 (
// Equation(s):
// \Selector12~7_combout  = (!ALUOp_EX[0] & (\portB~107_combout  & \Selector12~5_combout ))

	.dataa(gnd),
	.datab(ALUOp_EX_0),
	.datac(portB33),
	.datad(\Selector12~5_combout ),
	.cin(gnd),
	.combout(\Selector12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~7 .lut_mask = 16'h3000;
defparam \Selector12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N22
cycloneive_lcell_comb \Selector14~2 (
// Equation(s):
// \Selector14~2_combout  = (!\portB~103_combout  & (\ShiftLeft0~13_combout  & (!\ShiftLeft0~14_combout  & \Selector12~7_combout )))

	.dataa(portB32),
	.datab(\ShiftLeft0~13_combout ),
	.datac(\ShiftLeft0~14_combout ),
	.datad(\Selector12~7_combout ),
	.cin(gnd),
	.combout(\Selector14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~2 .lut_mask = 16'h0400;
defparam \Selector14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N24
cycloneive_lcell_comb \ShiftLeft0~64 (
// Equation(s):
// \ShiftLeft0~64_combout  = (\portB~92_combout  & (\portA~25_combout )) # (!\portB~92_combout  & ((\portA~67_combout )))

	.dataa(gnd),
	.datab(portA9),
	.datac(portA31),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~64 .lut_mask = 16'hCCF0;
defparam \ShiftLeft0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N22
cycloneive_lcell_comb \ShiftLeft0~65 (
// Equation(s):
// \ShiftLeft0~65_combout  = (\portB~97_combout  & (\ShiftLeft0~58_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~64_combout )))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftLeft0~58_combout ),
	.datad(\ShiftLeft0~64_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~65 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N16
cycloneive_lcell_comb \ShiftLeft0~66 (
// Equation(s):
// \ShiftLeft0~66_combout  = (\portB~100_combout  & ((\ShiftLeft0~53_combout ))) # (!\portB~100_combout  & (\ShiftLeft0~65_combout ))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftLeft0~65_combout ),
	.datad(\ShiftLeft0~53_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~66 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N0
cycloneive_lcell_comb \Selector12~8 (
// Equation(s):
// \Selector12~8_combout  = (ALUOp_EX[0]) # ((!\ShiftLeft0~16_combout  & ((\portB~103_combout ) # (\portB~107_combout ))))

	.dataa(ALUOp_EX_0),
	.datab(portB32),
	.datac(portB33),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~8 .lut_mask = 16'hAAFE;
defparam \Selector12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N22
cycloneive_lcell_comb \Selector12~9 (
// Equation(s):
// \Selector12~9_combout  = (\Selector12~5_combout  & !\Selector12~8_combout )

	.dataa(gnd),
	.datab(\Selector12~5_combout ),
	.datac(gnd),
	.datad(\Selector12~8_combout ),
	.cin(gnd),
	.combout(\Selector12~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~9 .lut_mask = 16'h00CC;
defparam \Selector12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N10
cycloneive_lcell_comb \Selector14~3 (
// Equation(s):
// \Selector14~3_combout  = (Selector12 & ((\ShiftRight0~29_combout ) # ((\ShiftLeft0~66_combout  & \Selector12~9_combout )))) # (!Selector12 & (\ShiftLeft0~66_combout  & (\Selector12~9_combout )))

	.dataa(Selector12),
	.datab(\ShiftLeft0~66_combout ),
	.datac(\Selector12~9_combout ),
	.datad(\ShiftRight0~29_combout ),
	.cin(gnd),
	.combout(\Selector14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~3 .lut_mask = 16'hEAC0;
defparam \Selector14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N4
cycloneive_lcell_comb \Selector14~4 (
// Equation(s):
// \Selector14~4_combout  = (\Selector14~1_combout ) # ((\Selector14~0_combout ) # ((\Selector14~2_combout ) # (\Selector14~3_combout )))

	.dataa(\Selector14~1_combout ),
	.datab(\Selector14~0_combout ),
	.datac(\Selector14~2_combout ),
	.datad(\Selector14~3_combout ),
	.cin(gnd),
	.combout(\Selector14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~4 .lut_mask = 16'hFFFE;
defparam \Selector14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N0
cycloneive_lcell_comb \Selector12~11 (
// Equation(s):
// \Selector12~11_combout  = (!ALUOp_EX[0] & (!\portB~107_combout  & (\portB~103_combout  & \Selector12~5_combout )))

	.dataa(ALUOp_EX_0),
	.datab(portB33),
	.datac(portB32),
	.datad(\Selector12~5_combout ),
	.cin(gnd),
	.combout(\Selector12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~11 .lut_mask = 16'h1000;
defparam \Selector12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N10
cycloneive_lcell_comb \Selector14~5 (
// Equation(s):
// \Selector14~5_combout  = (\Selector12~11_combout  & ((\portB~100_combout  & (\ShiftLeft0~23_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~39_combout )))))

	.dataa(portB31),
	.datab(\ShiftLeft0~23_combout ),
	.datac(\ShiftLeft0~39_combout ),
	.datad(\Selector12~11_combout ),
	.cin(gnd),
	.combout(\Selector14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~5 .lut_mask = 16'hD800;
defparam \Selector14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N0
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((\portB~62_combout  $ (\portA~25_combout  $ (\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((\portB~62_combout  & (\portA~25_combout  & !\Add1~31 )) # (!\portB~62_combout  & ((\portA~25_combout ) # (!\Add1~31 ))))

	.dataa(portB15),
	.datab(portA9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h964D;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N2
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (\portB~59_combout  & ((\portA~67_combout  & (!\Add1~33 )) # (!\portA~67_combout  & ((\Add1~33 ) # (GND))))) # (!\portB~59_combout  & ((\portA~67_combout  & (\Add1~33  & VCC)) # (!\portA~67_combout  & (!\Add1~33 ))))
// \Add1~35  = CARRY((\portB~59_combout  & ((!\Add1~33 ) # (!\portA~67_combout ))) # (!\portB~59_combout  & (!\portA~67_combout  & !\Add1~33 )))

	.dataa(portB14),
	.datab(portA31),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h692B;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N6
cycloneive_lcell_comb \Selector14~6 (
// Equation(s):
// \Selector14~6_combout  = (\Selector14~5_combout ) # ((\Selector0~11_combout  & \Add1~34_combout ))

	.dataa(\Selector0~11_combout ),
	.datab(gnd),
	.datac(\Selector14~5_combout ),
	.datad(\Add1~34_combout ),
	.cin(gnd),
	.combout(\Selector14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~6 .lut_mask = 16'hFAF0;
defparam \Selector14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N26
cycloneive_lcell_comb \Selector15~9 (
// Equation(s):
// \Selector15~9_combout  = (Selector12 & ((\portB~103_combout  & (\ShiftRight0~51_combout )) # (!\portB~103_combout  & ((\Selector23~0_combout )))))

	.dataa(Selector12),
	.datab(portB32),
	.datac(\ShiftRight0~51_combout ),
	.datad(\Selector23~0_combout ),
	.cin(gnd),
	.combout(\Selector15~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~9 .lut_mask = 16'hA280;
defparam \Selector15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N4
cycloneive_lcell_comb \Selector15~10 (
// Equation(s):
// \Selector15~10_combout  = (\Selector15~9_combout ) # ((\Selector0~11_combout  & \Add1~32_combout ))

	.dataa(\Selector15~9_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Add1~32_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~10 .lut_mask = 16'hEAEA;
defparam \Selector15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N20
cycloneive_lcell_comb \Selector15~5 (
// Equation(s):
// \Selector15~5_combout  = (\portB~62_combout  & (\Selector0~10_combout  & ((!\portA~25_combout )))) # (!\portB~62_combout  & ((\portA~25_combout  & (\Selector0~10_combout )) # (!\portA~25_combout  & ((\Selector0~13_combout )))))

	.dataa(portB15),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~13_combout ),
	.datad(portA9),
	.cin(gnd),
	.combout(\Selector15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~5 .lut_mask = 16'h44D8;
defparam \Selector15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N0
cycloneive_lcell_comb \Selector15~4 (
// Equation(s):
// \Selector15~4_combout  = (\portA~25_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \portB~62_combout )))) # (!\portA~25_combout  & (((\Selector0~8_combout  & \portB~62_combout ))))

	.dataa(\Selector0~9_combout ),
	.datab(portA9),
	.datac(\Selector0~8_combout ),
	.datad(portB15),
	.cin(gnd),
	.combout(\Selector15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~4 .lut_mask = 16'hF8C0;
defparam \Selector15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N14
cycloneive_lcell_comb \Selector15~6 (
// Equation(s):
// \Selector15~6_combout  = (\Selector12~11_combout  & ((\portB~100_combout  & ((\ShiftLeft0~28_combout ))) # (!\portB~100_combout  & (\ShiftLeft0~43_combout ))))

	.dataa(\ShiftLeft0~43_combout ),
	.datab(\ShiftLeft0~28_combout ),
	.datac(\Selector12~11_combout ),
	.datad(portB31),
	.cin(gnd),
	.combout(\Selector15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~6 .lut_mask = 16'hC0A0;
defparam \Selector15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N24
cycloneive_lcell_comb \ShiftLeft0~67 (
// Equation(s):
// \ShiftLeft0~67_combout  = (\portB~92_combout  & (\portA~27_combout )) # (!\portB~92_combout  & ((\portA~25_combout )))

	.dataa(portA10),
	.datab(portA9),
	.datac(gnd),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~67 .lut_mask = 16'hAACC;
defparam \ShiftLeft0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N26
cycloneive_lcell_comb \ShiftLeft0~68 (
// Equation(s):
// \ShiftLeft0~68_combout  = (\portB~97_combout  & (\ShiftLeft0~61_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~67_combout )))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftLeft0~61_combout ),
	.datad(\ShiftLeft0~67_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~68 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N2
cycloneive_lcell_comb \Selector15~12 (
// Equation(s):
// \Selector15~12_combout  = (\Selector12~9_combout  & ((\portB~100_combout  & (\ShiftLeft0~56_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~68_combout )))))

	.dataa(portB31),
	.datab(\ShiftLeft0~56_combout ),
	.datac(\ShiftLeft0~68_combout ),
	.datad(\Selector12~9_combout ),
	.cin(gnd),
	.combout(\Selector15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~12 .lut_mask = 16'hD800;
defparam \Selector15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N18
cycloneive_lcell_comb \Selector15~7 (
// Equation(s):
// \Selector15~7_combout  = (\Selector15~12_combout ) # ((!\ShiftLeft0~15_combout  & (\Selector12~7_combout  & \portA~69_combout )))

	.dataa(\ShiftLeft0~15_combout ),
	.datab(\Selector12~7_combout ),
	.datac(portA32),
	.datad(\Selector15~12_combout ),
	.cin(gnd),
	.combout(\Selector15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~7 .lut_mask = 16'hFF40;
defparam \Selector15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N12
cycloneive_lcell_comb \Selector15~8 (
// Equation(s):
// \Selector15~8_combout  = (\Selector15~5_combout ) # ((\Selector15~4_combout ) # ((\Selector15~6_combout ) # (\Selector15~7_combout )))

	.dataa(\Selector15~5_combout ),
	.datab(\Selector15~4_combout ),
	.datac(\Selector15~6_combout ),
	.datad(\Selector15~7_combout ),
	.cin(gnd),
	.combout(\Selector15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~8 .lut_mask = 16'hFFFE;
defparam \Selector15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N14
cycloneive_lcell_comb \Selector12~20 (
// Equation(s):
// \Selector12~20_combout  = (\ShiftLeft0~19_combout  & (!\portB~100_combout  & (!\portB~103_combout  & \Selector12~7_combout )))

	.dataa(\ShiftLeft0~19_combout ),
	.datab(portB31),
	.datac(portB32),
	.datad(\Selector12~7_combout ),
	.cin(gnd),
	.combout(\Selector12~20_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~20 .lut_mask = 16'h0200;
defparam \Selector12~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N4
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((\portA~65_combout  $ (\portB~56_combout  $ (\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((\portA~65_combout  & ((!\Add1~35 ) # (!\portB~56_combout ))) # (!\portA~65_combout  & (!\portB~56_combout  & !\Add1~35 )))

	.dataa(portA30),
	.datab(portB13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h962B;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N6
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (\portB~53_combout  & ((\portA~63_combout  & (!\Add1~37 )) # (!\portA~63_combout  & ((\Add1~37 ) # (GND))))) # (!\portB~53_combout  & ((\portA~63_combout  & (\Add1~37  & VCC)) # (!\portA~63_combout  & (!\Add1~37 ))))
// \Add1~39  = CARRY((\portB~53_combout  & ((!\Add1~37 ) # (!\portA~63_combout ))) # (!\portB~53_combout  & (!\portA~63_combout  & !\Add1~37 )))

	.dataa(portB12),
	.datab(portA29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h692B;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N28
cycloneive_lcell_comb \Selector12~17 (
// Equation(s):
// \Selector12~17_combout  = (\Selector12~20_combout ) # ((\Selector0~11_combout  & \Add1~38_combout ))

	.dataa(gnd),
	.datab(\Selector0~11_combout ),
	.datac(\Selector12~20_combout ),
	.datad(\Add1~38_combout ),
	.cin(gnd),
	.combout(\Selector12~17_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~17 .lut_mask = 16'hFCF0;
defparam \Selector12~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N4
cycloneive_lcell_comb \Add0~36 (
// Equation(s):
// \Add0~36_combout  = ((\portB~56_combout  $ (\portA~65_combout  $ (!\Add0~35 )))) # (GND)
// \Add0~37  = CARRY((\portB~56_combout  & ((\portA~65_combout ) # (!\Add0~35 ))) # (!\portB~56_combout  & (\portA~65_combout  & !\Add0~35 )))

	.dataa(portB13),
	.datab(portA30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~35 ),
	.combout(\Add0~36_combout ),
	.cout(\Add0~37 ));
// synopsys translate_off
defparam \Add0~36 .lut_mask = 16'h698E;
defparam \Add0~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N6
cycloneive_lcell_comb \Add0~38 (
// Equation(s):
// \Add0~38_combout  = (\portA~63_combout  & ((\portB~53_combout  & (\Add0~37  & VCC)) # (!\portB~53_combout  & (!\Add0~37 )))) # (!\portA~63_combout  & ((\portB~53_combout  & (!\Add0~37 )) # (!\portB~53_combout  & ((\Add0~37 ) # (GND)))))
// \Add0~39  = CARRY((\portA~63_combout  & (!\portB~53_combout  & !\Add0~37 )) # (!\portA~63_combout  & ((!\Add0~37 ) # (!\portB~53_combout ))))

	.dataa(portA29),
	.datab(portB12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~37 ),
	.combout(\Add0~38_combout ),
	.cout(\Add0~39 ));
// synopsys translate_off
defparam \Add0~38 .lut_mask = 16'h9617;
defparam \Add0~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N8
cycloneive_lcell_comb \Selector12~12 (
// Equation(s):
// \Selector12~12_combout  = (\portB~53_combout  & ((\Selector0~8_combout ) # ((\portA~63_combout  & \Selector0~9_combout )))) # (!\portB~53_combout  & (\portA~63_combout  & (\Selector0~8_combout )))

	.dataa(portB12),
	.datab(portA29),
	.datac(\Selector0~8_combout ),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~12 .lut_mask = 16'hE8E0;
defparam \Selector12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N22
cycloneive_lcell_comb \Selector12~13 (
// Equation(s):
// \Selector12~13_combout  = (\portA~63_combout  & (\Selector0~10_combout  & ((!\portB~53_combout )))) # (!\portA~63_combout  & ((\portB~53_combout  & (\Selector0~10_combout )) # (!\portB~53_combout  & ((\Selector0~13_combout )))))

	.dataa(portA29),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~13_combout ),
	.datad(portB12),
	.cin(gnd),
	.combout(\Selector12~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~13 .lut_mask = 16'h44D8;
defparam \Selector12~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N30
cycloneive_lcell_comb \Selector12~14 (
// Equation(s):
// \Selector12~14_combout  = (\Selector12~11_combout  & ((\portB~100_combout  & ((\ShiftLeft0~31_combout ))) # (!\portB~100_combout  & (\ShiftLeft0~45_combout ))))

	.dataa(\ShiftLeft0~45_combout ),
	.datab(\ShiftLeft0~31_combout ),
	.datac(portB31),
	.datad(\Selector12~11_combout ),
	.cin(gnd),
	.combout(\Selector12~14_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~14 .lut_mask = 16'hCA00;
defparam \Selector12~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N26
cycloneive_lcell_comb \ShiftLeft0~70 (
// Equation(s):
// \ShiftLeft0~70_combout  = (\portB~92_combout  & ((\portA~65_combout ))) # (!\portB~92_combout  & (\portA~63_combout ))

	.dataa(portA29),
	.datab(gnd),
	.datac(portA30),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~70 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N30
cycloneive_lcell_comb \ShiftLeft0~71 (
// Equation(s):
// \ShiftLeft0~71_combout  = (\portB~97_combout  & (\ShiftLeft0~64_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~70_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~64_combout ),
	.datac(portB30),
	.datad(\ShiftLeft0~70_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~71 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N0
cycloneive_lcell_comb \ShiftLeft0~72 (
// Equation(s):
// \ShiftLeft0~72_combout  = (\portB~100_combout  & (\ShiftLeft0~59_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~71_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~59_combout ),
	.datac(\ShiftLeft0~71_combout ),
	.datad(portB31),
	.cin(gnd),
	.combout(\ShiftLeft0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~72 .lut_mask = 16'hCCF0;
defparam \ShiftLeft0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N12
cycloneive_lcell_comb \Selector12~15 (
// Equation(s):
// \Selector12~15_combout  = (\Selector12~9_combout  & ((\ShiftLeft0~72_combout ) # ((Selector12 & \ShiftRight0~69_combout )))) # (!\Selector12~9_combout  & (((Selector12 & \ShiftRight0~69_combout ))))

	.dataa(\Selector12~9_combout ),
	.datab(\ShiftLeft0~72_combout ),
	.datac(Selector12),
	.datad(\ShiftRight0~69_combout ),
	.cin(gnd),
	.combout(\Selector12~15_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~15 .lut_mask = 16'hF888;
defparam \Selector12~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N18
cycloneive_lcell_comb \Selector12~16 (
// Equation(s):
// \Selector12~16_combout  = (\Selector12~12_combout ) # ((\Selector12~13_combout ) # ((\Selector12~14_combout ) # (\Selector12~15_combout )))

	.dataa(\Selector12~12_combout ),
	.datab(\Selector12~13_combout ),
	.datac(\Selector12~14_combout ),
	.datad(\Selector12~15_combout ),
	.cin(gnd),
	.combout(\Selector12~16_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~16 .lut_mask = 16'hFFFE;
defparam \Selector12~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N22
cycloneive_lcell_comb \Selector13~2 (
// Equation(s):
// \Selector13~2_combout  = (\portA~65_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & \portB~56_combout )))) # (!\portA~65_combout  & (((\Selector0~8_combout  & \portB~56_combout ))))

	.dataa(portA30),
	.datab(\Selector0~9_combout ),
	.datac(\Selector0~8_combout ),
	.datad(portB13),
	.cin(gnd),
	.combout(\Selector13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~2 .lut_mask = 16'hF8A0;
defparam \Selector13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N6
cycloneive_lcell_comb \Selector13~3 (
// Equation(s):
// \Selector13~3_combout  = (\portA~65_combout  & (((\Selector0~10_combout  & !\portB~56_combout )))) # (!\portA~65_combout  & ((\portB~56_combout  & ((\Selector0~10_combout ))) # (!\portB~56_combout  & (\Selector0~13_combout ))))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~10_combout ),
	.datac(portA30),
	.datad(portB13),
	.cin(gnd),
	.combout(\Selector13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~3 .lut_mask = 16'h0CCA;
defparam \Selector13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N14
cycloneive_lcell_comb \Selector13~4 (
// Equation(s):
// \Selector13~4_combout  = (\ShiftLeft0~75_combout  & ((\Selector12~9_combout ) # ((Selector12 & \ShiftRight0~78_combout )))) # (!\ShiftLeft0~75_combout  & (Selector12 & (\ShiftRight0~78_combout )))

	.dataa(\ShiftLeft0~75_combout ),
	.datab(Selector12),
	.datac(\ShiftRight0~78_combout ),
	.datad(\Selector12~9_combout ),
	.cin(gnd),
	.combout(\Selector13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~4 .lut_mask = 16'hEAC0;
defparam \Selector13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N16
cycloneive_lcell_comb \Selector13~9 (
// Equation(s):
// \Selector13~9_combout  = (!\portB~100_combout  & (\ShiftLeft0~21_combout  & (!\portB~103_combout  & \Selector12~7_combout )))

	.dataa(portB31),
	.datab(\ShiftLeft0~21_combout ),
	.datac(portB32),
	.datad(\Selector12~7_combout ),
	.cin(gnd),
	.combout(\Selector13~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~9 .lut_mask = 16'h0400;
defparam \Selector13~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N8
cycloneive_lcell_comb \Selector13~5 (
// Equation(s):
// \Selector13~5_combout  = (\Selector13~2_combout ) # ((\Selector13~3_combout ) # ((\Selector13~4_combout ) # (\Selector13~9_combout )))

	.dataa(\Selector13~2_combout ),
	.datab(\Selector13~3_combout ),
	.datac(\Selector13~4_combout ),
	.datad(\Selector13~9_combout ),
	.cin(gnd),
	.combout(\Selector13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~5 .lut_mask = 16'hFFFE;
defparam \Selector13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N20
cycloneive_lcell_comb \Selector13~6 (
// Equation(s):
// \Selector13~6_combout  = (\Selector12~11_combout  & ((\portB~100_combout  & ((\ShiftLeft0~34_combout ))) # (!\portB~100_combout  & (\ShiftLeft0~49_combout ))))

	.dataa(\ShiftLeft0~49_combout ),
	.datab(portB31),
	.datac(\ShiftLeft0~34_combout ),
	.datad(\Selector12~11_combout ),
	.cin(gnd),
	.combout(\Selector13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~6 .lut_mask = 16'hE200;
defparam \Selector13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N18
cycloneive_lcell_comb \Selector13~7 (
// Equation(s):
// \Selector13~7_combout  = (\Selector13~6_combout ) # ((\Selector0~11_combout  & \Add1~36_combout ))

	.dataa(\Selector0~11_combout ),
	.datab(gnd),
	.datac(\Add1~36_combout ),
	.datad(\Selector13~6_combout ),
	.cin(gnd),
	.combout(\Selector13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~7 .lut_mask = 16'hFFA0;
defparam \Selector13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N8
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = ((\portA~61_combout  $ (\portB~50_combout  $ (!\Add0~39 )))) # (GND)
// \Add0~41  = CARRY((\portA~61_combout  & ((\portB~50_combout ) # (!\Add0~39 ))) # (!\portA~61_combout  & (\portB~50_combout  & !\Add0~39 )))

	.dataa(portA28),
	.datab(portB11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~39 ),
	.combout(\Add0~40_combout ),
	.cout(\Add0~41 ));
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'h698E;
defparam \Add0~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N10
cycloneive_lcell_comb \Add0~42 (
// Equation(s):
// \Add0~42_combout  = (\portA~59_combout  & ((\portB~47_combout  & (\Add0~41  & VCC)) # (!\portB~47_combout  & (!\Add0~41 )))) # (!\portA~59_combout  & ((\portB~47_combout  & (!\Add0~41 )) # (!\portB~47_combout  & ((\Add0~41 ) # (GND)))))
// \Add0~43  = CARRY((\portA~59_combout  & (!\portB~47_combout  & !\Add0~41 )) # (!\portA~59_combout  & ((!\Add0~41 ) # (!\portB~47_combout ))))

	.dataa(portA27),
	.datab(portB10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~41 ),
	.combout(\Add0~42_combout ),
	.cout(\Add0~43 ));
// synopsys translate_off
defparam \Add0~42 .lut_mask = 16'h9617;
defparam \Add0~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N4
cycloneive_lcell_comb \Selector10~1 (
// Equation(s):
// \Selector10~1_combout  = (\Selector0~8_combout  & (((\portA~59_combout ) # (\portB~47_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\portA~59_combout  & \portB~47_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector0~8_combout ),
	.datac(portA27),
	.datad(portB10),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~1 .lut_mask = 16'hECC0;
defparam \Selector10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N14
cycloneive_lcell_comb \Selector10~2 (
// Equation(s):
// \Selector10~2_combout  = (\portA~59_combout  & (\Selector0~10_combout  & ((!\portB~47_combout )))) # (!\portA~59_combout  & ((\portB~47_combout  & (\Selector0~10_combout )) # (!\portB~47_combout  & ((\Selector0~13_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~13_combout ),
	.datac(portA27),
	.datad(portB10),
	.cin(gnd),
	.combout(\Selector10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~2 .lut_mask = 16'h0AAC;
defparam \Selector10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N30
cycloneive_lcell_comb \Selector10~3 (
// Equation(s):
// \Selector10~3_combout  = (\ShiftLeft0~24_combout  & (!\portB~103_combout  & \Selector12~7_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~24_combout ),
	.datac(portB32),
	.datad(\Selector12~7_combout ),
	.cin(gnd),
	.combout(\Selector10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~3 .lut_mask = 16'h0C00;
defparam \Selector10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N24
cycloneive_lcell_comb \Selector10~4 (
// Equation(s):
// \Selector10~4_combout  = (\ShiftLeft0~78_combout  & ((\Selector12~9_combout ) # ((Selector12 & \ShiftRight0~81_combout )))) # (!\ShiftLeft0~78_combout  & (Selector12 & ((\ShiftRight0~81_combout ))))

	.dataa(\ShiftLeft0~78_combout ),
	.datab(Selector12),
	.datac(\Selector12~9_combout ),
	.datad(\ShiftRight0~81_combout ),
	.cin(gnd),
	.combout(\Selector10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~4 .lut_mask = 16'hECA0;
defparam \Selector10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N22
cycloneive_lcell_comb \Selector10~5 (
// Equation(s):
// \Selector10~5_combout  = (\Selector10~1_combout ) # ((\Selector10~2_combout ) # ((\Selector10~3_combout ) # (\Selector10~4_combout )))

	.dataa(\Selector10~1_combout ),
	.datab(\Selector10~2_combout ),
	.datac(\Selector10~3_combout ),
	.datad(\Selector10~4_combout ),
	.cin(gnd),
	.combout(\Selector10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~5 .lut_mask = 16'hFFFE;
defparam \Selector10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N8
cycloneive_lcell_comb \Selector10~6 (
// Equation(s):
// \Selector10~6_combout  = (\Selector12~11_combout  & ((\portB~100_combout  & ((\ShiftLeft0~39_combout ))) # (!\portB~100_combout  & (\ShiftLeft0~53_combout ))))

	.dataa(\ShiftLeft0~53_combout ),
	.datab(portB31),
	.datac(\ShiftLeft0~39_combout ),
	.datad(\Selector12~11_combout ),
	.cin(gnd),
	.combout(\Selector10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~6 .lut_mask = 16'hE200;
defparam \Selector10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N8
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((\portB~50_combout  $ (\portA~61_combout  $ (\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((\portB~50_combout  & (\portA~61_combout  & !\Add1~39 )) # (!\portB~50_combout  & ((\portA~61_combout ) # (!\Add1~39 ))))

	.dataa(portB11),
	.datab(portA28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h964D;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N10
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (\portA~59_combout  & ((\portB~47_combout  & (!\Add1~41 )) # (!\portB~47_combout  & (\Add1~41  & VCC)))) # (!\portA~59_combout  & ((\portB~47_combout  & ((\Add1~41 ) # (GND))) # (!\portB~47_combout  & (!\Add1~41 ))))
// \Add1~43  = CARRY((\portA~59_combout  & (\portB~47_combout  & !\Add1~41 )) # (!\portA~59_combout  & ((\portB~47_combout ) # (!\Add1~41 ))))

	.dataa(portA27),
	.datab(portB10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h694D;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N2
cycloneive_lcell_comb \Selector10~7 (
// Equation(s):
// \Selector10~7_combout  = (\Selector10~6_combout ) # ((\Selector0~11_combout  & \Add1~42_combout ))

	.dataa(gnd),
	.datab(\Selector0~11_combout ),
	.datac(\Selector10~6_combout ),
	.datad(\Add1~42_combout ),
	.cin(gnd),
	.combout(\Selector10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~7 .lut_mask = 16'hFCF0;
defparam \Selector10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N24
cycloneive_lcell_comb \Selector11~2 (
// Equation(s):
// \Selector11~2_combout  = (\portA~61_combout  & (\Selector0~10_combout  & ((!\portB~50_combout )))) # (!\portA~61_combout  & ((\portB~50_combout  & (\Selector0~10_combout )) # (!\portB~50_combout  & ((\Selector0~13_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~13_combout ),
	.datac(portA28),
	.datad(portB11),
	.cin(gnd),
	.combout(\Selector11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~2 .lut_mask = 16'h0AAC;
defparam \Selector11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N4
cycloneive_lcell_comb \Selector11~1 (
// Equation(s):
// \Selector11~1_combout  = (\portA~61_combout  & ((\Selector0~8_combout ) # ((\portB~50_combout  & \Selector0~9_combout )))) # (!\portA~61_combout  & (\Selector0~8_combout  & (\portB~50_combout )))

	.dataa(portA28),
	.datab(\Selector0~8_combout ),
	.datac(portB11),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~1 .lut_mask = 16'hE8C8;
defparam \Selector11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N4
cycloneive_lcell_comb \Selector11~4 (
// Equation(s):
// \Selector11~4_combout  = (\ShiftLeft0~82_combout  & ((\Selector12~9_combout ) # ((\ShiftRight0~84_combout  & Selector12)))) # (!\ShiftLeft0~82_combout  & (\ShiftRight0~84_combout  & (Selector12)))

	.dataa(\ShiftLeft0~82_combout ),
	.datab(\ShiftRight0~84_combout ),
	.datac(Selector12),
	.datad(\Selector12~9_combout ),
	.cin(gnd),
	.combout(\Selector11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~4 .lut_mask = 16'hEAC0;
defparam \Selector11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N6
cycloneive_lcell_comb \Selector11~3 (
// Equation(s):
// \Selector11~3_combout  = (!\portB~103_combout  & (\ShiftLeft0~29_combout  & \Selector12~7_combout ))

	.dataa(gnd),
	.datab(portB32),
	.datac(\ShiftLeft0~29_combout ),
	.datad(\Selector12~7_combout ),
	.cin(gnd),
	.combout(\Selector11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~3 .lut_mask = 16'h3000;
defparam \Selector11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N30
cycloneive_lcell_comb \Selector11~5 (
// Equation(s):
// \Selector11~5_combout  = (\Selector11~2_combout ) # ((\Selector11~1_combout ) # ((\Selector11~4_combout ) # (\Selector11~3_combout )))

	.dataa(\Selector11~2_combout ),
	.datab(\Selector11~1_combout ),
	.datac(\Selector11~4_combout ),
	.datad(\Selector11~3_combout ),
	.cin(gnd),
	.combout(\Selector11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~5 .lut_mask = 16'hFFFE;
defparam \Selector11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N14
cycloneive_lcell_comb \Selector11~6 (
// Equation(s):
// \Selector11~6_combout  = (\Selector12~11_combout  & ((\portB~100_combout  & (\ShiftLeft0~43_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~56_combout )))))

	.dataa(portB31),
	.datab(\ShiftLeft0~43_combout ),
	.datac(\ShiftLeft0~56_combout ),
	.datad(\Selector12~11_combout ),
	.cin(gnd),
	.combout(\Selector11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~6 .lut_mask = 16'hD800;
defparam \Selector11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N28
cycloneive_lcell_comb \Selector11~7 (
// Equation(s):
// \Selector11~7_combout  = (\Selector11~6_combout ) # ((\Add1~40_combout  & \Selector0~11_combout ))

	.dataa(\Add1~40_combout ),
	.datab(\Selector0~11_combout ),
	.datac(gnd),
	.datad(\Selector11~6_combout ),
	.cin(gnd),
	.combout(\Selector11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~7 .lut_mask = 16'hFF88;
defparam \Selector11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N4
cycloneive_lcell_comb \Selector8~1 (
// Equation(s):
// \Selector8~1_combout  = (\portB~41_combout  & (((\Selector0~10_combout  & !\portA~55_combout )))) # (!\portB~41_combout  & ((\portA~55_combout  & ((\Selector0~10_combout ))) # (!\portA~55_combout  & (\Selector0~13_combout ))))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~10_combout ),
	.datac(portB8),
	.datad(portA25),
	.cin(gnd),
	.combout(\Selector8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~1 .lut_mask = 16'h0CCA;
defparam \Selector8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N2
cycloneive_lcell_comb \Selector8~5 (
// Equation(s):
// \Selector8~5_combout  = (\Selector0~8_combout  & (((\portB~41_combout ) # (\portA~55_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\portB~41_combout  & \portA~55_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(portB8),
	.datad(portA25),
	.cin(gnd),
	.combout(\Selector8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~5 .lut_mask = 16'hEAA0;
defparam \Selector8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N12
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((\portA~57_combout  $ (\portB~44_combout  $ (\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((\portA~57_combout  & ((!\Add1~43 ) # (!\portB~44_combout ))) # (!\portA~57_combout  & (!\portB~44_combout  & !\Add1~43 )))

	.dataa(portA26),
	.datab(portB9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h962B;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N14
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (\portA~55_combout  & ((\portB~41_combout  & (!\Add1~45 )) # (!\portB~41_combout  & (\Add1~45  & VCC)))) # (!\portA~55_combout  & ((\portB~41_combout  & ((\Add1~45 ) # (GND))) # (!\portB~41_combout  & (!\Add1~45 ))))
// \Add1~47  = CARRY((\portA~55_combout  & (\portB~41_combout  & !\Add1~45 )) # (!\portA~55_combout  & ((\portB~41_combout ) # (!\Add1~45 ))))

	.dataa(portA25),
	.datab(portB8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h694D;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N2
cycloneive_lcell_comb \Selector8~3 (
// Equation(s):
// \Selector8~3_combout  = (!\portB~103_combout  & (\ShiftLeft0~32_combout  & \Selector12~7_combout ))

	.dataa(portB32),
	.datab(gnd),
	.datac(\ShiftLeft0~32_combout ),
	.datad(\Selector12~7_combout ),
	.cin(gnd),
	.combout(\Selector8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~3 .lut_mask = 16'h5000;
defparam \Selector8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N24
cycloneive_lcell_comb \Selector8~4 (
// Equation(s):
// \Selector8~4_combout  = (\Selector8~2_combout ) # ((\Selector8~3_combout ) # ((\Selector8~0_combout  & \Selector12~11_combout )))

	.dataa(\Selector8~2_combout ),
	.datab(\Selector8~0_combout ),
	.datac(\Selector8~3_combout ),
	.datad(\Selector12~11_combout ),
	.cin(gnd),
	.combout(\Selector8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~4 .lut_mask = 16'hFEFA;
defparam \Selector8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N26
cycloneive_lcell_comb \Selector8~6 (
// Equation(s):
// \Selector8~6_combout  = (\Selector8~5_combout ) # ((\Selector8~4_combout ) # ((\Selector0~11_combout  & \Add1~46_combout )))

	.dataa(\Selector8~5_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Add1~46_combout ),
	.datad(\Selector8~4_combout ),
	.cin(gnd),
	.combout(\Selector8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~6 .lut_mask = 16'hFFEA;
defparam \Selector8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N12
cycloneive_lcell_comb \Add0~44 (
// Equation(s):
// \Add0~44_combout  = ((\portA~57_combout  $ (\portB~44_combout  $ (!\Add0~43 )))) # (GND)
// \Add0~45  = CARRY((\portA~57_combout  & ((\portB~44_combout ) # (!\Add0~43 ))) # (!\portA~57_combout  & (\portB~44_combout  & !\Add0~43 )))

	.dataa(portA26),
	.datab(portB9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~43 ),
	.combout(\Add0~44_combout ),
	.cout(\Add0~45 ));
// synopsys translate_off
defparam \Add0~44 .lut_mask = 16'h698E;
defparam \Add0~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N14
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// \Add0~46_combout  = (\portA~55_combout  & ((\portB~41_combout  & (\Add0~45  & VCC)) # (!\portB~41_combout  & (!\Add0~45 )))) # (!\portA~55_combout  & ((\portB~41_combout  & (!\Add0~45 )) # (!\portB~41_combout  & ((\Add0~45 ) # (GND)))))
// \Add0~47  = CARRY((\portA~55_combout  & (!\portB~41_combout  & !\Add0~45 )) # (!\portA~55_combout  & ((!\Add0~45 ) # (!\portB~41_combout ))))

	.dataa(portA25),
	.datab(portB8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~45 ),
	.combout(\Add0~46_combout ),
	.cout(\Add0~47 ));
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h9617;
defparam \Add0~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N14
cycloneive_lcell_comb \ShiftLeft0~85 (
// Equation(s):
// \ShiftLeft0~85_combout  = (\portB~92_combout  & (\portA~59_combout )) # (!\portB~92_combout  & ((\portA~57_combout )))

	.dataa(gnd),
	.datab(portA27),
	.datac(portB29),
	.datad(portA26),
	.cin(gnd),
	.combout(\ShiftLeft0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~85 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N20
cycloneive_lcell_comb \ShiftLeft0~80 (
// Equation(s):
// \ShiftLeft0~80_combout  = (\portB~92_combout  & (\portA~63_combout )) # (!\portB~92_combout  & ((\portA~61_combout )))

	.dataa(portA29),
	.datab(gnd),
	.datac(portA28),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~80 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N18
cycloneive_lcell_comb \ShiftLeft0~86 (
// Equation(s):
// \ShiftLeft0~86_combout  = (\portB~97_combout  & ((\ShiftLeft0~80_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~85_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftLeft0~85_combout ),
	.datad(\ShiftLeft0~80_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~86 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N26
cycloneive_lcell_comb \ShiftLeft0~74 (
// Equation(s):
// \ShiftLeft0~74_combout  = (!\portB~97_combout  & ((\portB~92_combout  & (\portA~67_combout )) # (!\portB~92_combout  & ((\portA~65_combout )))))

	.dataa(portB29),
	.datab(portA31),
	.datac(portB30),
	.datad(portA30),
	.cin(gnd),
	.combout(\ShiftLeft0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~74 .lut_mask = 16'h0D08;
defparam \ShiftLeft0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N16
cycloneive_lcell_comb \Selector1~0 (
// Equation(s):
// \Selector1~0_combout  = (\portB~100_combout  & ((\ShiftLeft0~73_combout ) # ((\ShiftLeft0~74_combout )))) # (!\portB~100_combout  & (((\ShiftLeft0~86_combout ))))

	.dataa(\ShiftLeft0~73_combout ),
	.datab(portB31),
	.datac(\ShiftLeft0~86_combout ),
	.datad(\ShiftLeft0~74_combout ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~0 .lut_mask = 16'hFCB8;
defparam \Selector1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N4
cycloneive_lcell_comb \Selector9~6 (
// Equation(s):
// \Selector9~6_combout  = (\Selector12~5_combout  & (!\Selector12~8_combout  & \Selector1~0_combout ))

	.dataa(\Selector12~5_combout ),
	.datab(gnd),
	.datac(\Selector12~8_combout ),
	.datad(\Selector1~0_combout ),
	.cin(gnd),
	.combout(\Selector9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~6 .lut_mask = 16'h0A00;
defparam \Selector9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N22
cycloneive_lcell_comb \Selector9~7 (
// Equation(s):
// \Selector9~7_combout  = (\Selector9~6_combout ) # ((\Selector0~11_combout  & \Add1~44_combout ))

	.dataa(gnd),
	.datab(\Selector0~11_combout ),
	.datac(\Selector9~6_combout ),
	.datad(\Add1~44_combout ),
	.cin(gnd),
	.combout(\Selector9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~7 .lut_mask = 16'hFCF0;
defparam \Selector9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N12
cycloneive_lcell_comb \Selector9~1 (
// Equation(s):
// \Selector9~1_combout  = (\portB~44_combout  & (\Selector0~10_combout  & (!\portA~57_combout ))) # (!\portB~44_combout  & ((\portA~57_combout  & (\Selector0~10_combout )) # (!\portA~57_combout  & ((\Selector0~13_combout )))))

	.dataa(portB9),
	.datab(\Selector0~10_combout ),
	.datac(portA26),
	.datad(\Selector0~13_combout ),
	.cin(gnd),
	.combout(\Selector9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~1 .lut_mask = 16'h4D48;
defparam \Selector9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N16
cycloneive_lcell_comb \Selector9~2 (
// Equation(s):
// \Selector9~2_combout  = (\Selector0~8_combout  & (((\portA~57_combout ) # (\portB~44_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\portA~57_combout  & \portB~44_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(portA26),
	.datad(portB9),
	.cin(gnd),
	.combout(\Selector9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~2 .lut_mask = 16'hEAA0;
defparam \Selector9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N4
cycloneive_lcell_comb \Selector9~3 (
// Equation(s):
// \Selector9~3_combout  = (!\portB~103_combout  & (\ShiftLeft0~35_combout  & \Selector12~7_combout ))

	.dataa(gnd),
	.datab(portB32),
	.datac(\ShiftLeft0~35_combout ),
	.datad(\Selector12~7_combout ),
	.cin(gnd),
	.combout(\Selector9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~3 .lut_mask = 16'h3000;
defparam \Selector9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N0
cycloneive_lcell_comb \Selector9~4 (
// Equation(s):
// \Selector9~4_combout  = (\Selector9~0_combout  & ((\Selector12~11_combout ) # ((Selector12 & \ShiftRight0~90_combout )))) # (!\Selector9~0_combout  & (Selector12 & (\ShiftRight0~90_combout )))

	.dataa(\Selector9~0_combout ),
	.datab(Selector12),
	.datac(\ShiftRight0~90_combout ),
	.datad(\Selector12~11_combout ),
	.cin(gnd),
	.combout(\Selector9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~4 .lut_mask = 16'hEAC0;
defparam \Selector9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N18
cycloneive_lcell_comb \Selector9~5 (
// Equation(s):
// \Selector9~5_combout  = (\Selector9~1_combout ) # ((\Selector9~2_combout ) # ((\Selector9~3_combout ) # (\Selector9~4_combout )))

	.dataa(\Selector9~1_combout ),
	.datab(\Selector9~2_combout ),
	.datac(\Selector9~3_combout ),
	.datad(\Selector9~4_combout ),
	.cin(gnd),
	.combout(\Selector9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~5 .lut_mask = 16'hFFFE;
defparam \Selector9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N16
cycloneive_lcell_comb \Add0~48 (
// Equation(s):
// \Add0~48_combout  = ((\portA~53_combout  $ (\portB~38_combout  $ (!\Add0~47 )))) # (GND)
// \Add0~49  = CARRY((\portA~53_combout  & ((\portB~38_combout ) # (!\Add0~47 ))) # (!\portA~53_combout  & (\portB~38_combout  & !\Add0~47 )))

	.dataa(portA24),
	.datab(portB7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~47 ),
	.combout(\Add0~48_combout ),
	.cout(\Add0~49 ));
// synopsys translate_off
defparam \Add0~48 .lut_mask = 16'h698E;
defparam \Add0~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N18
cycloneive_lcell_comb \Add0~50 (
// Equation(s):
// \Add0~50_combout  = (\portA~51_combout  & ((\portB~35_combout  & (\Add0~49  & VCC)) # (!\portB~35_combout  & (!\Add0~49 )))) # (!\portA~51_combout  & ((\portB~35_combout  & (!\Add0~49 )) # (!\portB~35_combout  & ((\Add0~49 ) # (GND)))))
// \Add0~51  = CARRY((\portA~51_combout  & (!\portB~35_combout  & !\Add0~49 )) # (!\portA~51_combout  & ((!\Add0~49 ) # (!\portB~35_combout ))))

	.dataa(portA23),
	.datab(portB6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~49 ),
	.combout(\Add0~50_combout ),
	.cout(\Add0~51 ));
// synopsys translate_off
defparam \Add0~50 .lut_mask = 16'h9617;
defparam \Add0~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N16
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((\portB~38_combout  $ (\portA~53_combout  $ (\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((\portB~38_combout  & (\portA~53_combout  & !\Add1~47 )) # (!\portB~38_combout  & ((\portA~53_combout ) # (!\Add1~47 ))))

	.dataa(portB7),
	.datab(portA24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h964D;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N18
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (\portA~51_combout  & ((\portB~35_combout  & (!\Add1~49 )) # (!\portB~35_combout  & (\Add1~49  & VCC)))) # (!\portA~51_combout  & ((\portB~35_combout  & ((\Add1~49 ) # (GND))) # (!\portB~35_combout  & (!\Add1~49 ))))
// \Add1~51  = CARRY((\portA~51_combout  & (\portB~35_combout  & !\Add1~49 )) # (!\portA~51_combout  & ((\portB~35_combout ) # (!\Add1~49 ))))

	.dataa(portA23),
	.datab(portB6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h694D;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N4
cycloneive_lcell_comb \Selector4~4 (
// Equation(s):
// \Selector4~4_combout  = (!\ShiftLeft0~7_combout  & (\Selector0~1_combout  & (!\ShiftLeft0~6_combout  & !\ShiftLeft0~10_combout )))

	.dataa(\ShiftLeft0~7_combout ),
	.datab(\Selector0~1_combout ),
	.datac(\ShiftLeft0~6_combout ),
	.datad(\ShiftLeft0~10_combout ),
	.cin(gnd),
	.combout(\Selector4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~4 .lut_mask = 16'h0004;
defparam \Selector4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N4
cycloneive_lcell_comb \ShiftLeft0~83 (
// Equation(s):
// \ShiftLeft0~83_combout  = (\portB~92_combout  & (\portA~57_combout )) # (!\portB~92_combout  & ((\portA~55_combout )))

	.dataa(gnd),
	.datab(portA26),
	.datac(portA25),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~83 .lut_mask = 16'hCCF0;
defparam \ShiftLeft0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N18
cycloneive_lcell_comb \ShiftLeft0~87 (
// Equation(s):
// \ShiftLeft0~87_combout  = (\portB~92_combout  & ((\portA~53_combout ))) # (!\portB~92_combout  & (\portA~51_combout ))

	.dataa(gnd),
	.datab(portA23),
	.datac(portA24),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~87 .lut_mask = 16'hF0CC;
defparam \ShiftLeft0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N20
cycloneive_lcell_comb \ShiftLeft0~88 (
// Equation(s):
// \ShiftLeft0~88_combout  = (\portB~97_combout  & (\ShiftLeft0~83_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~87_combout )))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftLeft0~83_combout ),
	.datad(\ShiftLeft0~87_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~88 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N14
cycloneive_lcell_comb \ShiftLeft0~76 (
// Equation(s):
// \ShiftLeft0~76_combout  = (\portB~92_combout  & ((\portA~61_combout ))) # (!\portB~92_combout  & (\portA~59_combout ))

	.dataa(gnd),
	.datab(portA27),
	.datac(portA28),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~76 .lut_mask = 16'hF0CC;
defparam \ShiftLeft0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N28
cycloneive_lcell_comb \ShiftLeft0~77 (
// Equation(s):
// \ShiftLeft0~77_combout  = (\portB~97_combout  & ((\ShiftLeft0~70_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~76_combout ))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftLeft0~76_combout ),
	.datad(\ShiftLeft0~70_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~77 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N22
cycloneive_lcell_comb \Selector6~1 (
// Equation(s):
// \Selector6~1_combout  = (\Selector4~0_combout  & ((\Selector4~1_combout ) # ((\ShiftLeft0~77_combout )))) # (!\Selector4~0_combout  & (!\Selector4~1_combout  & (\ShiftLeft0~88_combout )))

	.dataa(\Selector4~0_combout ),
	.datab(\Selector4~1_combout ),
	.datac(\ShiftLeft0~88_combout ),
	.datad(\ShiftLeft0~77_combout ),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~1 .lut_mask = 16'hBA98;
defparam \Selector6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N0
cycloneive_lcell_comb \Selector6~2 (
// Equation(s):
// \Selector6~2_combout  = (\Selector4~1_combout  & ((\Selector6~1_combout  & ((\ShiftLeft0~40_combout ))) # (!\Selector6~1_combout  & (\ShiftLeft0~66_combout )))) # (!\Selector4~1_combout  & (((\Selector6~1_combout ))))

	.dataa(\Selector4~1_combout ),
	.datab(\ShiftLeft0~66_combout ),
	.datac(\Selector6~1_combout ),
	.datad(\ShiftLeft0~40_combout ),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~2 .lut_mask = 16'hF858;
defparam \Selector6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N12
cycloneive_lcell_comb \Selector6~4 (
// Equation(s):
// \Selector6~4_combout  = (\Selector6~3_combout  & ((\Selector0~0_combout ) # ((\Selector4~4_combout  & \Selector6~2_combout )))) # (!\Selector6~3_combout  & (((\Selector4~4_combout  & \Selector6~2_combout ))))

	.dataa(\Selector6~3_combout ),
	.datab(\Selector0~0_combout ),
	.datac(\Selector4~4_combout ),
	.datad(\Selector6~2_combout ),
	.cin(gnd),
	.combout(\Selector6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~4 .lut_mask = 16'hF888;
defparam \Selector6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N18
cycloneive_lcell_comb \Selector6~6 (
// Equation(s):
// \Selector6~6_combout  = (Selector61) # ((\Selector6~4_combout ) # ((\Selector0~6_combout  & \Add1~50_combout )))

	.dataa(Selector61),
	.datab(\Selector0~6_combout ),
	.datac(\Add1~50_combout ),
	.datad(\Selector6~4_combout ),
	.cin(gnd),
	.combout(\Selector6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~6 .lut_mask = 16'hFFEA;
defparam \Selector6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N20
cycloneive_lcell_comb \Selector7~0 (
// Equation(s):
// \Selector7~0_combout  = (\portA~53_combout  & (((\Selector0~4_combout  & !\portB~38_combout )))) # (!\portA~53_combout  & ((\portB~38_combout  & ((\Selector0~4_combout ))) # (!\portB~38_combout  & (Selector0))))

	.dataa(Selector0),
	.datab(\Selector0~4_combout ),
	.datac(portA24),
	.datad(portB7),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~0 .lut_mask = 16'h0CCA;
defparam \Selector7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N14
cycloneive_lcell_comb \Selector7~1 (
// Equation(s):
// \Selector7~1_combout  = (\Selector0~0_combout  & (\ShiftRight0~51_combout  & !\Selector4~2_combout ))

	.dataa(\Selector0~0_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~51_combout ),
	.datad(\Selector4~2_combout ),
	.cin(gnd),
	.combout(\Selector7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~1 .lut_mask = 16'h00A0;
defparam \Selector7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N2
cycloneive_lcell_comb \ShiftLeft0~79 (
// Equation(s):
// \ShiftLeft0~79_combout  = (\portB~92_combout  & ((\portA~67_combout ))) # (!\portB~92_combout  & (\portA~65_combout ))

	.dataa(portA30),
	.datab(gnd),
	.datac(portA31),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~79 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N28
cycloneive_lcell_comb \ShiftLeft0~81 (
// Equation(s):
// \ShiftLeft0~81_combout  = (\portB~97_combout  & (\ShiftLeft0~79_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~80_combout )))

	.dataa(portB30),
	.datab(\ShiftLeft0~79_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~80_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~81 .lut_mask = 16'hDD88;
defparam \ShiftLeft0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N8
cycloneive_lcell_comb \ShiftLeft0~69 (
// Equation(s):
// \ShiftLeft0~69_combout  = (\portB~100_combout  & ((\ShiftLeft0~56_combout ))) # (!\portB~100_combout  & (\ShiftLeft0~68_combout ))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftLeft0~68_combout ),
	.datad(\ShiftLeft0~56_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~69 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N16
cycloneive_lcell_comb \ShiftLeft0~89 (
// Equation(s):
// \ShiftLeft0~89_combout  = (\portB~92_combout  & ((\portA~55_combout ))) # (!\portB~92_combout  & (\portA~53_combout ))

	.dataa(portA24),
	.datab(gnd),
	.datac(portB29),
	.datad(portA25),
	.cin(gnd),
	.combout(\ShiftLeft0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~89 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N30
cycloneive_lcell_comb \ShiftLeft0~90 (
// Equation(s):
// \ShiftLeft0~90_combout  = (\portB~97_combout  & (\ShiftLeft0~85_combout )) # (!\portB~97_combout  & ((\ShiftLeft0~89_combout )))

	.dataa(gnd),
	.datab(portB30),
	.datac(\ShiftLeft0~85_combout ),
	.datad(\ShiftLeft0~89_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~90 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N30
cycloneive_lcell_comb \Selector7~2 (
// Equation(s):
// \Selector7~2_combout  = (\Selector4~0_combout  & (((\Selector4~1_combout )))) # (!\Selector4~0_combout  & ((\Selector4~1_combout  & (\ShiftLeft0~69_combout )) # (!\Selector4~1_combout  & ((\ShiftLeft0~90_combout )))))

	.dataa(\Selector4~0_combout ),
	.datab(\ShiftLeft0~69_combout ),
	.datac(\ShiftLeft0~90_combout ),
	.datad(\Selector4~1_combout ),
	.cin(gnd),
	.combout(\Selector7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~2 .lut_mask = 16'hEE50;
defparam \Selector7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N24
cycloneive_lcell_comb \ShiftLeft0~97 (
// Equation(s):
// \ShiftLeft0~97_combout  = (\ShiftLeft0~41_combout ) # ((!\portB~100_combout  & (!\portB~103_combout  & \ShiftLeft0~43_combout )))

	.dataa(portB31),
	.datab(portB32),
	.datac(\ShiftLeft0~43_combout ),
	.datad(\ShiftLeft0~41_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~97 .lut_mask = 16'hFF10;
defparam \ShiftLeft0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N28
cycloneive_lcell_comb \Selector7~3 (
// Equation(s):
// \Selector7~3_combout  = (\Selector4~0_combout  & ((\Selector7~2_combout  & ((\ShiftLeft0~97_combout ))) # (!\Selector7~2_combout  & (\ShiftLeft0~81_combout )))) # (!\Selector4~0_combout  & (((\Selector7~2_combout ))))

	.dataa(\Selector4~0_combout ),
	.datab(\ShiftLeft0~81_combout ),
	.datac(\Selector7~2_combout ),
	.datad(\ShiftLeft0~97_combout ),
	.cin(gnd),
	.combout(\Selector7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~3 .lut_mask = 16'hF858;
defparam \Selector7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N8
cycloneive_lcell_comb \Selector7~4 (
// Equation(s):
// \Selector7~4_combout  = (\Selector7~0_combout ) # ((\Selector7~1_combout ) # ((\Selector4~4_combout  & \Selector7~3_combout )))

	.dataa(\Selector4~4_combout ),
	.datab(\Selector7~0_combout ),
	.datac(\Selector7~1_combout ),
	.datad(\Selector7~3_combout ),
	.cin(gnd),
	.combout(\Selector7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~4 .lut_mask = 16'hFEFC;
defparam \Selector7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N6
cycloneive_lcell_comb \Selector7~5 (
// Equation(s):
// \Selector7~5_combout  = (\Selector0~2_combout  & (((\portA~53_combout ) # (\portB~38_combout )))) # (!\Selector0~2_combout  & (\Selector0~3_combout  & (\portA~53_combout  & \portB~38_combout )))

	.dataa(\Selector0~3_combout ),
	.datab(\Selector0~2_combout ),
	.datac(portA24),
	.datad(portB7),
	.cin(gnd),
	.combout(\Selector7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~5 .lut_mask = 16'hECC0;
defparam \Selector7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N12
cycloneive_lcell_comb \Selector7~6 (
// Equation(s):
// \Selector7~6_combout  = (\Selector7~5_combout ) # ((\Selector0~6_combout  & \Add1~48_combout ))

	.dataa(\Selector7~5_combout ),
	.datab(gnd),
	.datac(\Selector0~6_combout ),
	.datad(\Add1~48_combout ),
	.cin(gnd),
	.combout(\Selector7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~6 .lut_mask = 16'hFAAA;
defparam \Selector7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N20
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// \Add0~52_combout  = ((\portB~32_combout  $ (\portA~49_combout  $ (!\Add0~51 )))) # (GND)
// \Add0~53  = CARRY((\portB~32_combout  & ((\portA~49_combout ) # (!\Add0~51 ))) # (!\portB~32_combout  & (\portA~49_combout  & !\Add0~51 )))

	.dataa(portB5),
	.datab(portA22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~51 ),
	.combout(\Add0~52_combout ),
	.cout(\Add0~53 ));
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'h698E;
defparam \Add0~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N22
cycloneive_lcell_comb \Add0~54 (
// Equation(s):
// \Add0~54_combout  = (\portA~47_combout  & ((\portB~29_combout  & (\Add0~53  & VCC)) # (!\portB~29_combout  & (!\Add0~53 )))) # (!\portA~47_combout  & ((\portB~29_combout  & (!\Add0~53 )) # (!\portB~29_combout  & ((\Add0~53 ) # (GND)))))
// \Add0~55  = CARRY((\portA~47_combout  & (!\portB~29_combout  & !\Add0~53 )) # (!\portA~47_combout  & ((!\Add0~53 ) # (!\portB~29_combout ))))

	.dataa(portA21),
	.datab(portB4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~53 ),
	.combout(\Add0~54_combout ),
	.cout(\Add0~55 ));
// synopsys translate_off
defparam \Add0~54 .lut_mask = 16'h9617;
defparam \Add0~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N18
cycloneive_lcell_comb \Selector4~10 (
// Equation(s):
// \Selector4~10_combout  = (\Selector0~2_combout  & ((\portA~47_combout ) # ((\portB~29_combout )))) # (!\Selector0~2_combout  & (\portA~47_combout  & (\Selector0~3_combout  & \portB~29_combout )))

	.dataa(\Selector0~2_combout ),
	.datab(portA21),
	.datac(\Selector0~3_combout ),
	.datad(portB4),
	.cin(gnd),
	.combout(\Selector4~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~10 .lut_mask = 16'hEA88;
defparam \Selector4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N20
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((\portA~49_combout  $ (\portB~32_combout  $ (\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((\portA~49_combout  & ((!\Add1~51 ) # (!\portB~32_combout ))) # (!\portA~49_combout  & (!\portB~32_combout  & !\Add1~51 )))

	.dataa(portA22),
	.datab(portB5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h962B;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N22
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (\portA~47_combout  & ((\portB~29_combout  & (!\Add1~53 )) # (!\portB~29_combout  & (\Add1~53  & VCC)))) # (!\portA~47_combout  & ((\portB~29_combout  & ((\Add1~53 ) # (GND))) # (!\portB~29_combout  & (!\Add1~53 ))))
// \Add1~55  = CARRY((\portA~47_combout  & (\portB~29_combout  & !\Add1~53 )) # (!\portA~47_combout  & ((\portB~29_combout ) # (!\Add1~53 ))))

	.dataa(portA21),
	.datab(portB4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h694D;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N30
cycloneive_lcell_comb \Selector4~11 (
// Equation(s):
// \Selector4~11_combout  = (\Selector4~10_combout ) # ((\Selector0~6_combout  & \Add1~54_combout ))

	.dataa(\Selector0~6_combout ),
	.datab(\Selector4~10_combout ),
	.datac(gnd),
	.datad(\Add1~54_combout ),
	.cin(gnd),
	.combout(\Selector4~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~11 .lut_mask = 16'hEECC;
defparam \Selector4~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N0
cycloneive_lcell_comb \Selector4~5 (
// Equation(s):
// \Selector4~5_combout  = (\portA~47_combout  & (((\Selector0~4_combout  & !\portB~29_combout )))) # (!\portA~47_combout  & ((\portB~29_combout  & ((\Selector0~4_combout ))) # (!\portB~29_combout  & (Selector0))))

	.dataa(Selector0),
	.datab(\Selector0~4_combout ),
	.datac(portA21),
	.datad(portB4),
	.cin(gnd),
	.combout(\Selector4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~5 .lut_mask = 16'h0CCA;
defparam \Selector4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N22
cycloneive_lcell_comb \Selector4~8 (
// Equation(s):
// \Selector4~8_combout  = (\Selector0~0_combout  & (\ShiftRight0~66_combout  & !\Selector4~2_combout ))

	.dataa(\Selector0~0_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~66_combout ),
	.datad(\Selector4~2_combout ),
	.cin(gnd),
	.combout(\Selector4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~8 .lut_mask = 16'h00A0;
defparam \Selector4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N14
cycloneive_lcell_comb \ShiftLeft0~84 (
// Equation(s):
// \ShiftLeft0~84_combout  = (\portB~97_combout  & ((\ShiftLeft0~76_combout ))) # (!\portB~97_combout  & (\ShiftLeft0~83_combout ))

	.dataa(portB30),
	.datab(gnd),
	.datac(\ShiftLeft0~83_combout ),
	.datad(\ShiftLeft0~76_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~84 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N26
cycloneive_lcell_comb \Selector4~6 (
// Equation(s):
// \Selector4~6_combout  = (\Selector4~1_combout  & (((\Selector4~0_combout )))) # (!\Selector4~1_combout  & ((\Selector4~0_combout  & ((\ShiftLeft0~84_combout ))) # (!\Selector4~0_combout  & (\ShiftLeft0~92_combout ))))

	.dataa(\ShiftLeft0~92_combout ),
	.datab(\Selector4~1_combout ),
	.datac(\Selector4~0_combout ),
	.datad(\ShiftLeft0~84_combout ),
	.cin(gnd),
	.combout(\Selector4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~6 .lut_mask = 16'hF2C2;
defparam \Selector4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N24
cycloneive_lcell_comb \Selector4~7 (
// Equation(s):
// \Selector4~7_combout  = (\Selector4~1_combout  & ((\Selector4~6_combout  & (\ShiftLeft0~47_combout )) # (!\Selector4~6_combout  & ((\ShiftLeft0~72_combout ))))) # (!\Selector4~1_combout  & (((\Selector4~6_combout ))))

	.dataa(\ShiftLeft0~47_combout ),
	.datab(\Selector4~1_combout ),
	.datac(\ShiftLeft0~72_combout ),
	.datad(\Selector4~6_combout ),
	.cin(gnd),
	.combout(\Selector4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~7 .lut_mask = 16'hBBC0;
defparam \Selector4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N20
cycloneive_lcell_comb \Selector4~9 (
// Equation(s):
// \Selector4~9_combout  = (\Selector4~5_combout ) # ((\Selector4~8_combout ) # ((\Selector4~4_combout  & \Selector4~7_combout )))

	.dataa(\Selector4~4_combout ),
	.datab(\Selector4~5_combout ),
	.datac(\Selector4~8_combout ),
	.datad(\Selector4~7_combout ),
	.cin(gnd),
	.combout(\Selector4~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~9 .lut_mask = 16'hFEFC;
defparam \Selector4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N28
cycloneive_lcell_comb \Selector5~0 (
// Equation(s):
// \Selector5~0_combout  = (\portB~32_combout  & (((\Selector0~4_combout  & !\portA~49_combout )))) # (!\portB~32_combout  & ((\portA~49_combout  & ((\Selector0~4_combout ))) # (!\portA~49_combout  & (Selector0))))

	.dataa(Selector0),
	.datab(\Selector0~4_combout ),
	.datac(portB5),
	.datad(portA22),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~0 .lut_mask = 16'h0CCA;
defparam \Selector5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N22
cycloneive_lcell_comb \Selector5~1 (
// Equation(s):
// \Selector5~1_combout  = (\Selector0~0_combout  & (\ShiftRight0~75_combout  & !\Selector4~2_combout ))

	.dataa(\Selector0~0_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~75_combout ),
	.datad(\Selector4~2_combout ),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~1 .lut_mask = 16'h00A0;
defparam \Selector5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N10
cycloneive_lcell_comb \ShiftLeft0~73 (
// Equation(s):
// \ShiftLeft0~73_combout  = (\portB~97_combout  & ((\portB~92_combout  & (\portA~27_combout )) # (!\portB~92_combout  & ((\portA~25_combout )))))

	.dataa(portA10),
	.datab(portB30),
	.datac(portB29),
	.datad(portA9),
	.cin(gnd),
	.combout(\ShiftLeft0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~73 .lut_mask = 16'h8C80;
defparam \ShiftLeft0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N24
cycloneive_lcell_comb \ShiftLeft0~75 (
// Equation(s):
// \ShiftLeft0~75_combout  = (\portB~100_combout  & (((\ShiftLeft0~62_combout )))) # (!\portB~100_combout  & ((\ShiftLeft0~73_combout ) # ((\ShiftLeft0~74_combout ))))

	.dataa(portB31),
	.datab(\ShiftLeft0~73_combout ),
	.datac(\ShiftLeft0~74_combout ),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~75 .lut_mask = 16'hFE54;
defparam \ShiftLeft0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N4
cycloneive_lcell_comb \Selector5~2 (
// Equation(s):
// \Selector5~2_combout  = (\Selector4~1_combout  & (((\Selector4~0_combout ) # (\ShiftLeft0~75_combout )))) # (!\Selector4~1_combout  & (\ShiftLeft0~94_combout  & (!\Selector4~0_combout )))

	.dataa(\ShiftLeft0~94_combout ),
	.datab(\Selector4~1_combout ),
	.datac(\Selector4~0_combout ),
	.datad(\ShiftLeft0~75_combout ),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~2 .lut_mask = 16'hCEC2;
defparam \Selector5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N18
cycloneive_lcell_comb \Selector5~3 (
// Equation(s):
// \Selector5~3_combout  = (\Selector4~0_combout  & ((\Selector5~2_combout  & ((\ShiftLeft0~51_combout ))) # (!\Selector5~2_combout  & (\ShiftLeft0~86_combout )))) # (!\Selector4~0_combout  & (((\Selector5~2_combout ))))

	.dataa(\ShiftLeft0~86_combout ),
	.datab(\Selector4~0_combout ),
	.datac(\Selector5~2_combout ),
	.datad(\ShiftLeft0~51_combout ),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~3 .lut_mask = 16'hF838;
defparam \Selector5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N24
cycloneive_lcell_comb \Selector5~4 (
// Equation(s):
// \Selector5~4_combout  = (\Selector5~0_combout ) # ((\Selector5~1_combout ) # ((\Selector4~4_combout  & \Selector5~3_combout )))

	.dataa(\Selector4~4_combout ),
	.datab(\Selector5~0_combout ),
	.datac(\Selector5~1_combout ),
	.datad(\Selector5~3_combout ),
	.cin(gnd),
	.combout(\Selector5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~4 .lut_mask = 16'hFEFC;
defparam \Selector5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N2
cycloneive_lcell_comb \Selector5~5 (
// Equation(s):
// \Selector5~5_combout  = (\Selector0~2_combout  & (((\portB~32_combout ) # (\portA~49_combout )))) # (!\Selector0~2_combout  & (\Selector0~3_combout  & (\portB~32_combout  & \portA~49_combout )))

	.dataa(\Selector0~3_combout ),
	.datab(\Selector0~2_combout ),
	.datac(portB5),
	.datad(portA22),
	.cin(gnd),
	.combout(\Selector5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~5 .lut_mask = 16'hECC0;
defparam \Selector5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N0
cycloneive_lcell_comb \Selector5~6 (
// Equation(s):
// \Selector5~6_combout  = (\Selector5~5_combout ) # ((\Selector0~6_combout  & \Add1~52_combout ))

	.dataa(\Selector0~6_combout ),
	.datab(gnd),
	.datac(\Selector5~5_combout ),
	.datad(\Add1~52_combout ),
	.cin(gnd),
	.combout(\Selector5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~6 .lut_mask = 16'hFAF0;
defparam \Selector5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N24
cycloneive_lcell_comb \Add0~56 (
// Equation(s):
// \Add0~56_combout  = ((\portA~45_combout  $ (\portB~26_combout  $ (!\Add0~55 )))) # (GND)
// \Add0~57  = CARRY((\portA~45_combout  & ((\portB~26_combout ) # (!\Add0~55 ))) # (!\portA~45_combout  & (\portB~26_combout  & !\Add0~55 )))

	.dataa(portA20),
	.datab(portB3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~55 ),
	.combout(\Add0~56_combout ),
	.cout(\Add0~57 ));
// synopsys translate_off
defparam \Add0~56 .lut_mask = 16'h698E;
defparam \Add0~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N26
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// \Add0~58_combout  = (\portA~41_combout  & ((\portB~23_combout  & (\Add0~57  & VCC)) # (!\portB~23_combout  & (!\Add0~57 )))) # (!\portA~41_combout  & ((\portB~23_combout  & (!\Add0~57 )) # (!\portB~23_combout  & ((\Add0~57 ) # (GND)))))
// \Add0~59  = CARRY((\portA~41_combout  & (!\portB~23_combout  & !\Add0~57 )) # (!\portA~41_combout  & ((!\Add0~57 ) # (!\portB~23_combout ))))

	.dataa(portA18),
	.datab(portB2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~57 ),
	.combout(\Add0~58_combout ),
	.cout(\Add0~59 ));
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'h9617;
defparam \Add0~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N28
cycloneive_lcell_comb \Selector2~3 (
// Equation(s):
// \Selector2~3_combout  = (\Selector0~8_combout  & (((\portA~41_combout ) # (\portB~23_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\portA~41_combout  & \portB~23_combout )))

	.dataa(\Selector0~9_combout ),
	.datab(\Selector0~8_combout ),
	.datac(portA18),
	.datad(portB2),
	.cin(gnd),
	.combout(\Selector2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~3 .lut_mask = 16'hECC0;
defparam \Selector2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N24
cycloneive_lcell_comb \Selector2~9 (
// Equation(s):
// \Selector2~9_combout  = (\portA~41_combout  & (\Selector0~10_combout  & ((!\portB~23_combout )))) # (!\portA~41_combout  & ((\portB~23_combout  & (\Selector0~10_combout )) # (!\portB~23_combout  & ((\Selector0~13_combout )))))

	.dataa(\Selector0~10_combout ),
	.datab(\Selector0~13_combout ),
	.datac(portA18),
	.datad(portB2),
	.cin(gnd),
	.combout(\Selector2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~9 .lut_mask = 16'h0AAC;
defparam \Selector2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N10
cycloneive_lcell_comb \ShiftLeft0~78 (
// Equation(s):
// \ShiftLeft0~78_combout  = (\portB~100_combout  & (\ShiftLeft0~65_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~77_combout )))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftLeft0~65_combout ),
	.datad(\ShiftLeft0~77_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~78 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N28
cycloneive_lcell_comb \Selector2~4 (
// Equation(s):
// \Selector2~4_combout  = (\ShiftLeft0~17_combout  & (\ShiftLeft0~95_combout  & (!\Selector2~2_combout ))) # (!\ShiftLeft0~17_combout  & (((\Selector2~2_combout ) # (\ShiftLeft0~88_combout ))))

	.dataa(\ShiftLeft0~95_combout ),
	.datab(\ShiftLeft0~17_combout ),
	.datac(\Selector2~2_combout ),
	.datad(\ShiftLeft0~88_combout ),
	.cin(gnd),
	.combout(\Selector2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~4 .lut_mask = 16'h3B38;
defparam \Selector2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N26
cycloneive_lcell_comb \Selector2~5 (
// Equation(s):
// \Selector2~5_combout  = (\Selector2~2_combout  & ((\Selector2~4_combout  & ((\ShiftLeft0~78_combout ))) # (!\Selector2~4_combout  & (\ShiftLeft0~91_combout )))) # (!\Selector2~2_combout  & (((\Selector2~4_combout ))))

	.dataa(\ShiftLeft0~91_combout ),
	.datab(\ShiftLeft0~78_combout ),
	.datac(\Selector2~2_combout ),
	.datad(\Selector2~4_combout ),
	.cin(gnd),
	.combout(\Selector2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~5 .lut_mask = 16'hCFA0;
defparam \Selector2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N12
cycloneive_lcell_comb \Selector2~6 (
// Equation(s):
// \Selector2~6_combout  = (ALUOp_EX[0]) # ((ALUOp_EX[1]) # ((\portB~107_combout  & !\ShiftLeft0~16_combout )))

	.dataa(portB33),
	.datab(ALUOp_EX_0),
	.datac(ALUOp_EX_1),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~6 .lut_mask = 16'hFCFE;
defparam \Selector2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N22
cycloneive_lcell_comb \Selector2~7 (
// Equation(s):
// \Selector2~7_combout  = (\Selector12~19_combout  & (\Selector2~5_combout  & !\Selector2~6_combout ))

	.dataa(gnd),
	.datab(\Selector12~19_combout ),
	.datac(\Selector2~5_combout ),
	.datad(\Selector2~6_combout ),
	.cin(gnd),
	.combout(\Selector2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~7 .lut_mask = 16'h00C0;
defparam \Selector2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N26
cycloneive_lcell_comb \Selector2~12 (
// Equation(s):
// \Selector2~12_combout  = (!\portB~100_combout  & (\ShiftRight0~18_combout  & (!\portB~103_combout  & Selector12)))

	.dataa(portB31),
	.datab(\ShiftRight0~18_combout ),
	.datac(portB32),
	.datad(Selector12),
	.cin(gnd),
	.combout(\Selector2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~12 .lut_mask = 16'h0400;
defparam \Selector2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N8
cycloneive_lcell_comb \Selector2~8 (
// Equation(s):
// \Selector2~8_combout  = (\Selector2~7_combout ) # ((\Selector2~12_combout ) # ((\ShiftLeft0~54_combout  & \Selector12~7_combout )))

	.dataa(\ShiftLeft0~54_combout ),
	.datab(\Selector12~7_combout ),
	.datac(\Selector2~7_combout ),
	.datad(\Selector2~12_combout ),
	.cin(gnd),
	.combout(\Selector2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~8 .lut_mask = 16'hFFF8;
defparam \Selector2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N24
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((\portA~45_combout  $ (\portB~26_combout  $ (\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((\portA~45_combout  & ((!\Add1~55 ) # (!\portB~26_combout ))) # (!\portA~45_combout  & (!\portB~26_combout  & !\Add1~55 )))

	.dataa(portA20),
	.datab(portB3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h962B;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N26
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = (\portB~23_combout  & ((\portA~41_combout  & (!\Add1~57 )) # (!\portA~41_combout  & ((\Add1~57 ) # (GND))))) # (!\portB~23_combout  & ((\portA~41_combout  & (\Add1~57  & VCC)) # (!\portA~41_combout  & (!\Add1~57 ))))
// \Add1~59  = CARRY((\portB~23_combout  & ((!\Add1~57 ) # (!\portA~41_combout ))) # (!\portB~23_combout  & (!\portA~41_combout  & !\Add1~57 )))

	.dataa(portB2),
	.datab(portA18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout(\Add1~59 ));
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'h692B;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N10
cycloneive_lcell_comb \Selector2~10 (
// Equation(s):
// \Selector2~10_combout  = (\Selector2~9_combout ) # ((\Selector2~8_combout ) # ((\Selector0~11_combout  & \Add1~58_combout )))

	.dataa(\Selector2~9_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Selector2~8_combout ),
	.datad(\Add1~58_combout ),
	.cin(gnd),
	.combout(\Selector2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~10 .lut_mask = 16'hFEFA;
defparam \Selector2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N18
cycloneive_lcell_comb \Selector3~2 (
// Equation(s):
// \Selector3~2_combout  = (\portA~45_combout  & ((\Selector0~8_combout ) # ((\portB~26_combout  & \Selector0~9_combout )))) # (!\portA~45_combout  & (\Selector0~8_combout  & (\portB~26_combout )))

	.dataa(portA20),
	.datab(\Selector0~8_combout ),
	.datac(portB3),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~2 .lut_mask = 16'hE8C8;
defparam \Selector3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N12
cycloneive_lcell_comb \Selector3~7 (
// Equation(s):
// \Selector3~7_combout  = (\portA~45_combout  & (((\Selector0~10_combout  & !\portB~26_combout )))) # (!\portA~45_combout  & ((\portB~26_combout  & ((\Selector0~10_combout ))) # (!\portB~26_combout  & (\Selector0~13_combout ))))

	.dataa(portA20),
	.datab(\Selector0~13_combout ),
	.datac(\Selector0~10_combout ),
	.datad(portB3),
	.cin(gnd),
	.combout(\Selector3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~7 .lut_mask = 16'h50E4;
defparam \Selector3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N10
cycloneive_lcell_comb \Selector3~10 (
// Equation(s):
// \Selector3~10_combout  = (!\portB~100_combout  & (!\portB~103_combout  & (\ShiftRight0~47_combout  & Selector12)))

	.dataa(portB31),
	.datab(portB32),
	.datac(\ShiftRight0~47_combout ),
	.datad(Selector12),
	.cin(gnd),
	.combout(\Selector3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~10 .lut_mask = 16'h1000;
defparam \Selector3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N20
cycloneive_lcell_comb \ShiftLeft0~93 (
// Equation(s):
// \ShiftLeft0~93_combout  = (\portB~92_combout  & ((\portA~51_combout ))) # (!\portB~92_combout  & (\portA~49_combout ))

	.dataa(gnd),
	.datab(portA22),
	.datac(portB29),
	.datad(portA23),
	.cin(gnd),
	.combout(\ShiftLeft0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~93 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N8
cycloneive_lcell_comb \ShiftLeft0~96 (
// Equation(s):
// \ShiftLeft0~96_combout  = (\portB~92_combout  & ((\portA~47_combout ))) # (!\portB~92_combout  & (\portA~45_combout ))

	.dataa(gnd),
	.datab(portB29),
	.datac(portA20),
	.datad(portA21),
	.cin(gnd),
	.combout(\ShiftLeft0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~96 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N30
cycloneive_lcell_comb \Selector3~3 (
// Equation(s):
// \Selector3~3_combout  = (\Selector2~2_combout  & (((!\ShiftLeft0~17_combout )))) # (!\Selector2~2_combout  & ((\ShiftLeft0~17_combout  & ((\ShiftLeft0~96_combout ))) # (!\ShiftLeft0~17_combout  & (\ShiftLeft0~90_combout ))))

	.dataa(\Selector2~2_combout ),
	.datab(\ShiftLeft0~90_combout ),
	.datac(\ShiftLeft0~17_combout ),
	.datad(\ShiftLeft0~96_combout ),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~3 .lut_mask = 16'h5E0E;
defparam \Selector3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N16
cycloneive_lcell_comb \ShiftLeft0~82 (
// Equation(s):
// \ShiftLeft0~82_combout  = (\portB~100_combout  & (\ShiftLeft0~68_combout )) # (!\portB~100_combout  & ((\ShiftLeft0~81_combout )))

	.dataa(gnd),
	.datab(portB31),
	.datac(\ShiftLeft0~68_combout ),
	.datad(\ShiftLeft0~81_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~82 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N0
cycloneive_lcell_comb \Selector3~4 (
// Equation(s):
// \Selector3~4_combout  = (\Selector2~2_combout  & ((\Selector3~3_combout  & ((\ShiftLeft0~82_combout ))) # (!\Selector3~3_combout  & (\ShiftLeft0~93_combout )))) # (!\Selector2~2_combout  & (((\Selector3~3_combout ))))

	.dataa(\Selector2~2_combout ),
	.datab(\ShiftLeft0~93_combout ),
	.datac(\Selector3~3_combout ),
	.datad(\ShiftLeft0~82_combout ),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~4 .lut_mask = 16'hF858;
defparam \Selector3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N2
cycloneive_lcell_comb \Selector3~5 (
// Equation(s):
// \Selector3~5_combout  = (\Selector3~4_combout  & (\Selector12~19_combout  & !\Selector2~6_combout ))

	.dataa(gnd),
	.datab(\Selector3~4_combout ),
	.datac(\Selector12~19_combout ),
	.datad(\Selector2~6_combout ),
	.cin(gnd),
	.combout(\Selector3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~5 .lut_mask = 16'h00C0;
defparam \Selector3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N4
cycloneive_lcell_comb \Selector3~6 (
// Equation(s):
// \Selector3~6_combout  = (\Selector3~10_combout ) # ((\Selector3~5_combout ) # ((ShiftLeft0 & \Selector12~7_combout )))

	.dataa(ShiftLeft0),
	.datab(\Selector12~7_combout ),
	.datac(\Selector3~10_combout ),
	.datad(\Selector3~5_combout ),
	.cin(gnd),
	.combout(\Selector3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~6 .lut_mask = 16'hFFF8;
defparam \Selector3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N18
cycloneive_lcell_comb \Selector3~8 (
// Equation(s):
// \Selector3~8_combout  = (\Selector3~7_combout ) # ((\Selector3~6_combout ) # ((\Selector0~11_combout  & \Add1~56_combout )))

	.dataa(\Selector0~11_combout ),
	.datab(\Selector3~7_combout ),
	.datac(\Selector3~6_combout ),
	.datad(\Add1~56_combout ),
	.cin(gnd),
	.combout(\Selector3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~8 .lut_mask = 16'hFEFC;
defparam \Selector3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N28
cycloneive_lcell_comb \Add0~60 (
// Equation(s):
// \Add0~60_combout  = ((\portA~43_combout  $ (\portB~20_combout  $ (!\Add0~59 )))) # (GND)
// \Add0~61  = CARRY((\portA~43_combout  & ((\portB~20_combout ) # (!\Add0~59 ))) # (!\portA~43_combout  & (\portB~20_combout  & !\Add0~59 )))

	.dataa(portA19),
	.datab(portB1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~59 ),
	.combout(\Add0~60_combout ),
	.cout(\Add0~61 ));
// synopsys translate_off
defparam \Add0~60 .lut_mask = 16'h698E;
defparam \Add0~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N30
cycloneive_lcell_comb \Add0~62 (
// Equation(s):
// \Add0~62_combout  = \portA~39_combout  $ (\Add0~61  $ (\portB~17_combout ))

	.dataa(portA17),
	.datab(gnd),
	.datac(gnd),
	.datad(portB),
	.cin(\Add0~61 ),
	.combout(\Add0~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~62 .lut_mask = 16'hA55A;
defparam \Add0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N14
cycloneive_lcell_comb \Selector0~17 (
// Equation(s):
// \Selector0~17_combout  = (\portB~17_combout  & ((\Selector0~8_combout ) # ((\Selector0~10_combout  & !\portA~39_combout )))) # (!\portB~17_combout  & (((\Selector0~10_combout  & \portA~39_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~10_combout ),
	.datac(portA17),
	.datad(portB),
	.cin(gnd),
	.combout(\Selector0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~17 .lut_mask = 16'hAEC0;
defparam \Selector0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N0
cycloneive_lcell_comb \Selector0~18 (
// Equation(s):
// \Selector0~18_combout  = (\Selector0~8_combout ) # ((\Selector0~9_combout  & \portB~17_combout ))

	.dataa(\Selector0~8_combout ),
	.datab(gnd),
	.datac(\Selector0~9_combout ),
	.datad(portB),
	.cin(gnd),
	.combout(\Selector0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~18 .lut_mask = 16'hFAAA;
defparam \Selector0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N22
cycloneive_lcell_comb \Selector0~19 (
// Equation(s):
// \Selector0~19_combout  = (\portA~39_combout  & ((\Selector0~18_combout ) # ((Selector12 & !\ShiftLeft0~15_combout ))))

	.dataa(portA17),
	.datab(Selector12),
	.datac(\ShiftLeft0~15_combout ),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~19 .lut_mask = 16'hAA08;
defparam \Selector0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N28
cycloneive_lcell_comb \Add1~60 (
// Equation(s):
// \Add1~60_combout  = ((\portB~20_combout  $ (\portA~43_combout  $ (\Add1~59 )))) # (GND)
// \Add1~61  = CARRY((\portB~20_combout  & (\portA~43_combout  & !\Add1~59 )) # (!\portB~20_combout  & ((\portA~43_combout ) # (!\Add1~59 ))))

	.dataa(portB1),
	.datab(portA19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~59 ),
	.combout(\Add1~60_combout ),
	.cout(\Add1~61 ));
// synopsys translate_off
defparam \Add1~60 .lut_mask = 16'h964D;
defparam \Add1~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N30
cycloneive_lcell_comb \Add1~62 (
// Equation(s):
// \Add1~62_combout  = \portB~17_combout  $ (\Add1~61  $ (!\portA~39_combout ))

	.dataa(gnd),
	.datab(portB),
	.datac(gnd),
	.datad(portA17),
	.cin(\Add1~61 ),
	.combout(\Add1~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~62 .lut_mask = 16'h3CC3;
defparam \Add1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N8
cycloneive_lcell_comb \Selector0~20 (
// Equation(s):
// \Selector0~20_combout  = (\Selector0~13_combout  & (!\portA~39_combout  & !\portB~17_combout ))

	.dataa(gnd),
	.datab(\Selector0~13_combout ),
	.datac(portA17),
	.datad(portB),
	.cin(gnd),
	.combout(\Selector0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~20 .lut_mask = 16'h000C;
defparam \Selector0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N30
cycloneive_lcell_comb \Selector0~21 (
// Equation(s):
// \Selector0~21_combout  = (\portB~100_combout ) # ((\portB~92_combout  & !\portB~97_combout ))

	.dataa(gnd),
	.datab(portB29),
	.datac(portB30),
	.datad(portB31),
	.cin(gnd),
	.combout(\Selector0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~21 .lut_mask = 16'hFF0C;
defparam \Selector0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N10
cycloneive_lcell_comb \ShiftLeft0~95 (
// Equation(s):
// \ShiftLeft0~95_combout  = (\portB~92_combout  & (\portA~45_combout )) # (!\portB~92_combout  & ((\portA~41_combout )))

	.dataa(portA20),
	.datab(gnd),
	.datac(portA18),
	.datad(portB29),
	.cin(gnd),
	.combout(\ShiftLeft0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~95 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N2
cycloneive_lcell_comb \Selector0~22 (
// Equation(s):
// \Selector0~22_combout  = (\ShiftLeft0~14_combout  & (((\Selector0~21_combout ) # (\ShiftLeft0~95_combout )))) # (!\ShiftLeft0~14_combout  & (\portA~39_combout  & (!\Selector0~21_combout )))

	.dataa(portA17),
	.datab(\ShiftLeft0~14_combout ),
	.datac(\Selector0~21_combout ),
	.datad(\ShiftLeft0~95_combout ),
	.cin(gnd),
	.combout(\Selector0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~22 .lut_mask = 16'hCEC2;
defparam \Selector0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N20
cycloneive_lcell_comb \Selector0~23 (
// Equation(s):
// \Selector0~23_combout  = (\Selector0~21_combout  & ((\Selector0~22_combout  & (\ShiftLeft0~92_combout )) # (!\Selector0~22_combout  & ((\portA~43_combout ))))) # (!\Selector0~21_combout  & (((\Selector0~22_combout ))))

	.dataa(\ShiftLeft0~92_combout ),
	.datab(portA19),
	.datac(\Selector0~21_combout ),
	.datad(\Selector0~22_combout ),
	.cin(gnd),
	.combout(\Selector0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~23 .lut_mask = 16'hAFC0;
defparam \Selector0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N18
cycloneive_lcell_comb \Selector0~24 (
// Equation(s):
// \Selector0~24_combout  = (\Selector12~9_combout  & ((\Selector0~23_combout ) # ((\Selector12~7_combout  & \ShiftLeft0~60_combout )))) # (!\Selector12~9_combout  & (((\Selector12~7_combout  & \ShiftLeft0~60_combout ))))

	.dataa(\Selector12~9_combout ),
	.datab(\Selector0~23_combout ),
	.datac(\Selector12~7_combout ),
	.datad(\ShiftLeft0~60_combout ),
	.cin(gnd),
	.combout(\Selector0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~24 .lut_mask = 16'hF888;
defparam \Selector0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N28
cycloneive_lcell_comb \Selector0~25 (
// Equation(s):
// \Selector0~25_combout  = (\Selector0~20_combout ) # ((\Selector0~24_combout ) # ((\Selector0~16_combout  & \Selector12~11_combout )))

	.dataa(\Selector0~16_combout ),
	.datab(\Selector12~11_combout ),
	.datac(\Selector0~20_combout ),
	.datad(\Selector0~24_combout ),
	.cin(gnd),
	.combout(\Selector0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~25 .lut_mask = 16'hFFF8;
defparam \Selector0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N10
cycloneive_lcell_comb \Selector0~26 (
// Equation(s):
// \Selector0~26_combout  = (\Selector0~19_combout ) # ((\Selector0~25_combout ) # ((\Selector0~11_combout  & \Add1~62_combout )))

	.dataa(\Selector0~19_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Add1~62_combout ),
	.datad(\Selector0~25_combout ),
	.cin(gnd),
	.combout(\Selector0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~26 .lut_mask = 16'hFFEA;
defparam \Selector0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N20
cycloneive_lcell_comb \Selector1~1 (
// Equation(s):
// \Selector1~1_combout  = (\ShiftRight0~45_combout  & (!\ShiftLeft0~14_combout  & (Selector12 & !\portB~103_combout )))

	.dataa(\ShiftRight0~45_combout ),
	.datab(\ShiftLeft0~14_combout ),
	.datac(Selector12),
	.datad(portB32),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~1 .lut_mask = 16'h0020;
defparam \Selector1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N0
cycloneive_lcell_comb \Selector1~7 (
// Equation(s):
// \Selector1~7_combout  = (\Selector0~8_combout  & (((\portA~43_combout ) # (\portB~20_combout )))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\portA~43_combout  & \portB~20_combout )))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(portA19),
	.datad(portB1),
	.cin(gnd),
	.combout(\Selector1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~7 .lut_mask = 16'hEAA0;
defparam \Selector1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N12
cycloneive_lcell_comb \Selector1~5 (
// Equation(s):
// \Selector1~5_combout  = (\Selector1~4_combout  & ((\Selector12~9_combout ) # ((\Selector12~7_combout  & \ShiftLeft0~63_combout )))) # (!\Selector1~4_combout  & (\Selector12~7_combout  & (\ShiftLeft0~63_combout )))

	.dataa(\Selector1~4_combout ),
	.datab(\Selector12~7_combout ),
	.datac(\ShiftLeft0~63_combout ),
	.datad(\Selector12~9_combout ),
	.cin(gnd),
	.combout(\Selector1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~5 .lut_mask = 16'hEAC0;
defparam \Selector1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N22
cycloneive_lcell_comb \Selector1~6 (
// Equation(s):
// \Selector1~6_combout  = (\Selector1~2_combout ) # ((\Selector1~5_combout ) # ((\Selector1~0_combout  & \Selector12~11_combout )))

	.dataa(\Selector1~2_combout ),
	.datab(\Selector1~0_combout ),
	.datac(\Selector12~11_combout ),
	.datad(\Selector1~5_combout ),
	.cin(gnd),
	.combout(\Selector1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~6 .lut_mask = 16'hFFEA;
defparam \Selector1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N0
cycloneive_lcell_comb \Selector1~8 (
// Equation(s):
// \Selector1~8_combout  = (\Selector1~7_combout ) # ((\Selector1~6_combout ) # ((\Selector0~11_combout  & \Add1~60_combout )))

	.dataa(\Selector1~7_combout ),
	.datab(\Selector0~11_combout ),
	.datac(\Selector1~6_combout ),
	.datad(\Add1~60_combout ),
	.cin(gnd),
	.combout(\Selector1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~8 .lut_mask = 16'hFEFA;
defparam \Selector1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N30
cycloneive_lcell_comb \Selector7~8 (
// Equation(s):
// \Selector7~8_combout  = (!\portB~107_combout  & (\Selector0~0_combout  & (!\portB~103_combout  & !\ShiftLeft0~16_combout )))

	.dataa(portB33),
	.datab(\Selector0~0_combout ),
	.datac(portB32),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\Selector7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~8 .lut_mask = 16'h0004;
defparam \Selector7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N4
cycloneive_lcell_comb \Selector31~6 (
// Equation(s):
// \Selector31~6_combout  = (Selector0 & (!\portA~69_combout  & !\portB~92_combout ))

	.dataa(gnd),
	.datab(Selector0),
	.datac(portA32),
	.datad(portB29),
	.cin(gnd),
	.combout(\Selector31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~6 .lut_mask = 16'h000C;
defparam \Selector31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N2
cycloneive_lcell_comb \ShiftRight0~86 (
// Equation(s):
// \ShiftRight0~86_combout  = (\portB~100_combout  & (((!\portB~103_combout  & \ShiftRight0~65_combout )))) # (!\portB~100_combout  & (\ShiftRight0~63_combout  & (\portB~103_combout )))

	.dataa(portB31),
	.datab(\ShiftRight0~63_combout ),
	.datac(portB32),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~86 .lut_mask = 16'h4A40;
defparam \ShiftRight0~86 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module btb (
	pc_out_3,
	pc_out_2,
	pc_out_5,
	pc_out_4,
	pc_out_7,
	pc_out_6,
	pc_out_9,
	pc_out_8,
	pc_out_11,
	pc_out_10,
	pc_out_13,
	pc_out_12,
	pc_out_15,
	pc_out_14,
	pc_out_17,
	pc_out_16,
	pc_out_19,
	pc_out_18,
	pc_out_21,
	pc_out_20,
	pc_out_23,
	pc_out_22,
	pc_out_25,
	pc_out_24,
	pc_out_27,
	pc_out_26,
	pc_out_29,
	pc_out_28,
	pc_out_31,
	pc_out_30,
	btbframesframeblocks2tag_1,
	btbframesframeblocks1tag_1,
	btbframesframeblocks0tag_1,
	btbframesframeblocks3tag_1,
	btbframesframeblocks1tag_0,
	btbframesframeblocks2tag_0,
	btbframesframeblocks0tag_0,
	btbframesframeblocks3tag_0,
	btbframesframeblocks2tag_3,
	btbframesframeblocks1tag_3,
	btbframesframeblocks0tag_3,
	btbframesframeblocks3tag_3,
	btbframesframeblocks1tag_2,
	btbframesframeblocks2tag_2,
	btbframesframeblocks0tag_2,
	btbframesframeblocks3tag_2,
	btbframesframeblocks2tag_5,
	btbframesframeblocks1tag_5,
	btbframesframeblocks0tag_5,
	btbframesframeblocks3tag_5,
	btbframesframeblocks1tag_4,
	btbframesframeblocks2tag_4,
	btbframesframeblocks0tag_4,
	btbframesframeblocks3tag_4,
	btbframesframeblocks2tag_7,
	btbframesframeblocks1tag_7,
	btbframesframeblocks0tag_7,
	btbframesframeblocks3tag_7,
	btbframesframeblocks1tag_6,
	btbframesframeblocks2tag_6,
	btbframesframeblocks0tag_6,
	btbframesframeblocks3tag_6,
	btbframesframeblocks2tag_9,
	btbframesframeblocks1tag_9,
	btbframesframeblocks0tag_9,
	btbframesframeblocks3tag_9,
	btbframesframeblocks1tag_8,
	btbframesframeblocks2tag_8,
	btbframesframeblocks0tag_8,
	btbframesframeblocks3tag_8,
	btbframesframeblocks2tag_11,
	btbframesframeblocks1tag_11,
	btbframesframeblocks0tag_11,
	btbframesframeblocks3tag_11,
	btbframesframeblocks1tag_10,
	btbframesframeblocks2tag_10,
	btbframesframeblocks0tag_10,
	btbframesframeblocks3tag_10,
	btbframesframeblocks2tag_13,
	btbframesframeblocks1tag_13,
	btbframesframeblocks0tag_13,
	btbframesframeblocks3tag_13,
	btbframesframeblocks1tag_12,
	btbframesframeblocks2tag_12,
	btbframesframeblocks0tag_12,
	btbframesframeblocks3tag_12,
	btbframesframeblocks2tag_15,
	btbframesframeblocks1tag_15,
	btbframesframeblocks0tag_15,
	btbframesframeblocks3tag_15,
	btbframesframeblocks1tag_14,
	btbframesframeblocks2tag_14,
	btbframesframeblocks0tag_14,
	btbframesframeblocks3tag_14,
	btbframesframeblocks2tag_17,
	btbframesframeblocks1tag_17,
	btbframesframeblocks0tag_17,
	btbframesframeblocks3tag_17,
	btbframesframeblocks1tag_16,
	btbframesframeblocks2tag_16,
	btbframesframeblocks0tag_16,
	btbframesframeblocks3tag_16,
	btbframesframeblocks2tag_19,
	btbframesframeblocks1tag_19,
	btbframesframeblocks0tag_19,
	btbframesframeblocks3tag_19,
	btbframesframeblocks1tag_18,
	btbframesframeblocks2tag_18,
	btbframesframeblocks0tag_18,
	btbframesframeblocks3tag_18,
	btbframesframeblocks2tag_21,
	btbframesframeblocks1tag_21,
	btbframesframeblocks0tag_21,
	btbframesframeblocks3tag_21,
	btbframesframeblocks1tag_20,
	btbframesframeblocks2tag_20,
	btbframesframeblocks0tag_20,
	btbframesframeblocks3tag_20,
	btbframesframeblocks2tag_23,
	btbframesframeblocks1tag_23,
	btbframesframeblocks0tag_23,
	btbframesframeblocks3tag_23,
	btbframesframeblocks1tag_22,
	btbframesframeblocks2tag_22,
	btbframesframeblocks0tag_22,
	btbframesframeblocks3tag_22,
	btbframesframeblocks2tag_25,
	btbframesframeblocks1tag_25,
	btbframesframeblocks0tag_25,
	btbframesframeblocks3tag_25,
	btbframesframeblocks1tag_24,
	btbframesframeblocks2tag_24,
	btbframesframeblocks0tag_24,
	btbframesframeblocks3tag_24,
	btbframesframeblocks2tag_27,
	btbframesframeblocks1tag_27,
	btbframesframeblocks0tag_27,
	btbframesframeblocks3tag_27,
	btbframesframeblocks1tag_26,
	btbframesframeblocks2tag_26,
	btbframesframeblocks0tag_26,
	btbframesframeblocks3tag_26,
	btbframesframeblocks2valid,
	btbframesframeblocks1valid,
	btbframesframeblocks0valid,
	btbframesframeblocks3valid,
	btbframesframeblocks1curr_state_1,
	btbframesframeblocks2curr_state_1,
	btbframesframeblocks0curr_state_1,
	btbframesframeblocks3curr_state_1,
	predicted,
	devpor,
	devclrn,
	devoe);
input 	pc_out_3;
input 	pc_out_2;
input 	pc_out_5;
input 	pc_out_4;
input 	pc_out_7;
input 	pc_out_6;
input 	pc_out_9;
input 	pc_out_8;
input 	pc_out_11;
input 	pc_out_10;
input 	pc_out_13;
input 	pc_out_12;
input 	pc_out_15;
input 	pc_out_14;
input 	pc_out_17;
input 	pc_out_16;
input 	pc_out_19;
input 	pc_out_18;
input 	pc_out_21;
input 	pc_out_20;
input 	pc_out_23;
input 	pc_out_22;
input 	pc_out_25;
input 	pc_out_24;
input 	pc_out_27;
input 	pc_out_26;
input 	pc_out_29;
input 	pc_out_28;
input 	pc_out_31;
input 	pc_out_30;
input 	btbframesframeblocks2tag_1;
input 	btbframesframeblocks1tag_1;
input 	btbframesframeblocks0tag_1;
input 	btbframesframeblocks3tag_1;
input 	btbframesframeblocks1tag_0;
input 	btbframesframeblocks2tag_0;
input 	btbframesframeblocks0tag_0;
input 	btbframesframeblocks3tag_0;
input 	btbframesframeblocks2tag_3;
input 	btbframesframeblocks1tag_3;
input 	btbframesframeblocks0tag_3;
input 	btbframesframeblocks3tag_3;
input 	btbframesframeblocks1tag_2;
input 	btbframesframeblocks2tag_2;
input 	btbframesframeblocks0tag_2;
input 	btbframesframeblocks3tag_2;
input 	btbframesframeblocks2tag_5;
input 	btbframesframeblocks1tag_5;
input 	btbframesframeblocks0tag_5;
input 	btbframesframeblocks3tag_5;
input 	btbframesframeblocks1tag_4;
input 	btbframesframeblocks2tag_4;
input 	btbframesframeblocks0tag_4;
input 	btbframesframeblocks3tag_4;
input 	btbframesframeblocks2tag_7;
input 	btbframesframeblocks1tag_7;
input 	btbframesframeblocks0tag_7;
input 	btbframesframeblocks3tag_7;
input 	btbframesframeblocks1tag_6;
input 	btbframesframeblocks2tag_6;
input 	btbframesframeblocks0tag_6;
input 	btbframesframeblocks3tag_6;
input 	btbframesframeblocks2tag_9;
input 	btbframesframeblocks1tag_9;
input 	btbframesframeblocks0tag_9;
input 	btbframesframeblocks3tag_9;
input 	btbframesframeblocks1tag_8;
input 	btbframesframeblocks2tag_8;
input 	btbframesframeblocks0tag_8;
input 	btbframesframeblocks3tag_8;
input 	btbframesframeblocks2tag_11;
input 	btbframesframeblocks1tag_11;
input 	btbframesframeblocks0tag_11;
input 	btbframesframeblocks3tag_11;
input 	btbframesframeblocks1tag_10;
input 	btbframesframeblocks2tag_10;
input 	btbframesframeblocks0tag_10;
input 	btbframesframeblocks3tag_10;
input 	btbframesframeblocks2tag_13;
input 	btbframesframeblocks1tag_13;
input 	btbframesframeblocks0tag_13;
input 	btbframesframeblocks3tag_13;
input 	btbframesframeblocks1tag_12;
input 	btbframesframeblocks2tag_12;
input 	btbframesframeblocks0tag_12;
input 	btbframesframeblocks3tag_12;
input 	btbframesframeblocks2tag_15;
input 	btbframesframeblocks1tag_15;
input 	btbframesframeblocks0tag_15;
input 	btbframesframeblocks3tag_15;
input 	btbframesframeblocks1tag_14;
input 	btbframesframeblocks2tag_14;
input 	btbframesframeblocks0tag_14;
input 	btbframesframeblocks3tag_14;
input 	btbframesframeblocks2tag_17;
input 	btbframesframeblocks1tag_17;
input 	btbframesframeblocks0tag_17;
input 	btbframesframeblocks3tag_17;
input 	btbframesframeblocks1tag_16;
input 	btbframesframeblocks2tag_16;
input 	btbframesframeblocks0tag_16;
input 	btbframesframeblocks3tag_16;
input 	btbframesframeblocks2tag_19;
input 	btbframesframeblocks1tag_19;
input 	btbframesframeblocks0tag_19;
input 	btbframesframeblocks3tag_19;
input 	btbframesframeblocks1tag_18;
input 	btbframesframeblocks2tag_18;
input 	btbframesframeblocks0tag_18;
input 	btbframesframeblocks3tag_18;
input 	btbframesframeblocks2tag_21;
input 	btbframesframeblocks1tag_21;
input 	btbframesframeblocks0tag_21;
input 	btbframesframeblocks3tag_21;
input 	btbframesframeblocks1tag_20;
input 	btbframesframeblocks2tag_20;
input 	btbframesframeblocks0tag_20;
input 	btbframesframeblocks3tag_20;
input 	btbframesframeblocks2tag_23;
input 	btbframesframeblocks1tag_23;
input 	btbframesframeblocks0tag_23;
input 	btbframesframeblocks3tag_23;
input 	btbframesframeblocks1tag_22;
input 	btbframesframeblocks2tag_22;
input 	btbframesframeblocks0tag_22;
input 	btbframesframeblocks3tag_22;
input 	btbframesframeblocks2tag_25;
input 	btbframesframeblocks1tag_25;
input 	btbframesframeblocks0tag_25;
input 	btbframesframeblocks3tag_25;
input 	btbframesframeblocks1tag_24;
input 	btbframesframeblocks2tag_24;
input 	btbframesframeblocks0tag_24;
input 	btbframesframeblocks3tag_24;
input 	btbframesframeblocks2tag_27;
input 	btbframesframeblocks1tag_27;
input 	btbframesframeblocks0tag_27;
input 	btbframesframeblocks3tag_27;
input 	btbframesframeblocks1tag_26;
input 	btbframesframeblocks2tag_26;
input 	btbframesframeblocks0tag_26;
input 	btbframesframeblocks3tag_26;
input 	btbframesframeblocks2valid;
input 	btbframesframeblocks1valid;
input 	btbframesframeblocks0valid;
input 	btbframesframeblocks3valid;
input 	btbframesframeblocks1curr_state_1;
input 	btbframesframeblocks2curr_state_1;
input 	btbframesframeblocks0curr_state_1;
input 	btbframesframeblocks3curr_state_1;
output 	predicted;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux21~0_combout ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \Mux16~0_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux12~0_combout ;
wire \Mux7~0_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux4~0_combout ;
wire \Mux1~0_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux4~1_combout ;
wire \predicted~15_combout ;
wire \Mux1~1_combout ;
wire \predicted~16_combout ;
wire \predicted~17_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \predicted~11_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \predicted~13_combout ;
wire \Mux7~1_combout ;
wire \predicted~12_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Mux12~1_combout ;
wire \predicted~10_combout ;
wire \predicted~14_combout ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \predicted~5_combout ;
wire \Mux16~1_combout ;
wire \predicted~7_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \predicted~6_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \predicted~8_combout ;
wire \predicted~9_combout ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \predicted~0_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \predicted~2_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \Mux21~1_combout ;
wire \predicted~3_combout ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \predicted~1_combout ;
wire \predicted~4_combout ;


// Location: LCCOMB_X53_Y40_N12
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].tag [3])) # (!pc_out_2 & ((\btbframes.frameblocks[0].tag [3])))))

	.dataa(btbframesframeblocks1tag_3),
	.datab(pc_out_3),
	.datac(pc_out_2),
	.datad(btbframesframeblocks0tag_3),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hE3E0;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N16
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\Mux25~0_combout  & (((\btbframes.frameblocks[3].tag [3])) # (!pc_out_3))) # (!\Mux25~0_combout  & (pc_out_3 & (\btbframes.frameblocks[2].tag [3])))

	.dataa(\Mux25~0_combout ),
	.datab(pc_out_3),
	.datac(btbframesframeblocks2tag_3),
	.datad(btbframesframeblocks3tag_3),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hEA62;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N0
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (pc_out_3 & (pc_out_2)) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].tag [7])) # (!pc_out_2 & ((\btbframes.frameblocks[0].tag [7])))))

	.dataa(pc_out_3),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_7),
	.datad(btbframesframeblocks0tag_7),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hD9C8;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N20
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (pc_out_2 & (pc_out_3)) # (!pc_out_2 & ((pc_out_3 & (\btbframes.frameblocks[2].tag [8])) # (!pc_out_3 & ((\btbframes.frameblocks[0].tag [8])))))

	.dataa(pc_out_2),
	.datab(pc_out_3),
	.datac(btbframesframeblocks2tag_8),
	.datad(btbframesframeblocks0tag_8),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hD9C8;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N26
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (\Mux20~0_combout  & (((\btbframes.frameblocks[3].tag [8])) # (!pc_out_2))) # (!\Mux20~0_combout  & (pc_out_2 & (\btbframes.frameblocks[1].tag [8])))

	.dataa(\Mux20~0_combout ),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_8),
	.datad(btbframesframeblocks3tag_8),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hEA62;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N14
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (pc_out_2 & (pc_out_3)) # (!pc_out_2 & ((pc_out_3 & (\btbframes.frameblocks[2].tag [10])) # (!pc_out_3 & ((\btbframes.frameblocks[0].tag [10])))))

	.dataa(pc_out_2),
	.datab(pc_out_3),
	.datac(btbframesframeblocks2tag_10),
	.datad(btbframesframeblocks0tag_10),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hD9C8;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N12
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (pc_out_2 & ((\Mux18~0_combout  & ((\btbframes.frameblocks[3].tag [10]))) # (!\Mux18~0_combout  & (\btbframes.frameblocks[1].tag [10])))) # (!pc_out_2 & (\Mux18~0_combout ))

	.dataa(pc_out_2),
	.datab(\Mux18~0_combout ),
	.datac(btbframesframeblocks1tag_10),
	.datad(btbframesframeblocks3tag_10),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hEC64;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N14
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (pc_out_2 & (((\btbframes.frameblocks[1].tag [13]) # (pc_out_3)))) # (!pc_out_2 & (\btbframes.frameblocks[0].tag [13] & ((!pc_out_3))))

	.dataa(btbframesframeblocks0tag_13),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_13),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hCCE2;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N20
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (\Mux15~0_combout  & (((\btbframes.frameblocks[3].tag [13])) # (!pc_out_3))) # (!\Mux15~0_combout  & (pc_out_3 & ((\btbframes.frameblocks[2].tag [13]))))

	.dataa(\Mux15~0_combout ),
	.datab(pc_out_3),
	.datac(btbframesframeblocks3tag_13),
	.datad(btbframesframeblocks2tag_13),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hE6A2;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N22
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (pc_out_2 & (((pc_out_3)))) # (!pc_out_2 & ((pc_out_3 & ((\btbframes.frameblocks[2].tag [12]))) # (!pc_out_3 & (\btbframes.frameblocks[0].tag [12]))))

	.dataa(pc_out_2),
	.datab(btbframesframeblocks0tag_12),
	.datac(btbframesframeblocks2tag_12),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hFA44;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N20
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (pc_out_2 & (((\btbframes.frameblocks[1].tag [15]) # (pc_out_3)))) # (!pc_out_2 & (\btbframes.frameblocks[0].tag [15] & ((!pc_out_3))))

	.dataa(btbframesframeblocks0tag_15),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_15),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hCCE2;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N14
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (pc_out_3 & ((\Mux13~0_combout  & (\btbframes.frameblocks[3].tag [15])) # (!\Mux13~0_combout  & ((\btbframes.frameblocks[2].tag [15]))))) # (!pc_out_3 & (((\Mux13~0_combout ))))

	.dataa(btbframesframeblocks3tag_15),
	.datab(pc_out_3),
	.datac(btbframesframeblocks2tag_15),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hBBC0;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N6
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (pc_out_2 & (((pc_out_3)))) # (!pc_out_2 & ((pc_out_3 & (\btbframes.frameblocks[2].tag [16])) # (!pc_out_3 & ((\btbframes.frameblocks[0].tag [16])))))

	.dataa(btbframesframeblocks2tag_16),
	.datab(pc_out_2),
	.datac(pc_out_3),
	.datad(btbframesframeblocks0tag_16),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hE3E0;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N30
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & ((\btbframes.frameblocks[1].tag [21]))) # (!pc_out_2 & (\btbframes.frameblocks[0].tag [21]))))

	.dataa(btbframesframeblocks0tag_21),
	.datab(pc_out_3),
	.datac(btbframesframeblocks1tag_21),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hFC22;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N6
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (pc_out_2 & (((pc_out_3)))) # (!pc_out_2 & ((pc_out_3 & (\btbframes.frameblocks[2].tag [20])) # (!pc_out_3 & ((\btbframes.frameblocks[0].tag [20])))))

	.dataa(pc_out_2),
	.datab(btbframesframeblocks2tag_20),
	.datac(btbframesframeblocks0tag_20),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hEE50;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N26
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (pc_out_2 & ((\Mux8~0_combout  & (\btbframes.frameblocks[3].tag [20])) # (!\Mux8~0_combout  & ((\btbframes.frameblocks[1].tag [20]))))) # (!pc_out_2 & (((\Mux8~0_combout ))))

	.dataa(btbframesframeblocks3tag_20),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_20),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hBBC0;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N12
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].tag [23])) # (!pc_out_2 & ((\btbframes.frameblocks[0].tag [23])))))

	.dataa(pc_out_3),
	.datab(btbframesframeblocks1tag_23),
	.datac(btbframesframeblocks0tag_23),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hEE50;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N14
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (pc_out_3 & ((\Mux5~0_combout  & ((\btbframes.frameblocks[3].tag [23]))) # (!\Mux5~0_combout  & (\btbframes.frameblocks[2].tag [23])))) # (!pc_out_3 & (((\Mux5~0_combout ))))

	.dataa(pc_out_3),
	.datab(btbframesframeblocks2tag_23),
	.datac(btbframesframeblocks3tag_23),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hF588;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N24
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (pc_out_2 & (((\btbframes.frameblocks[1].tag [25]) # (pc_out_3)))) # (!pc_out_2 & (\btbframes.frameblocks[0].tag [25] & ((!pc_out_3))))

	.dataa(btbframesframeblocks0tag_25),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_25),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hCCE2;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N22
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (\Mux3~0_combout  & (((\btbframes.frameblocks[3].tag [25])) # (!pc_out_3))) # (!\Mux3~0_combout  & (pc_out_3 & ((\btbframes.frameblocks[2].tag [25]))))

	.dataa(\Mux3~0_combout ),
	.datab(pc_out_3),
	.datac(btbframesframeblocks3tag_25),
	.datad(btbframesframeblocks2tag_25),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hE6A2;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N8
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (pc_out_3 & (((\btbframes.frameblocks[2].tag [24]) # (pc_out_2)))) # (!pc_out_3 & (\btbframes.frameblocks[0].tag [24] & ((!pc_out_2))))

	.dataa(btbframesframeblocks0tag_24),
	.datab(pc_out_3),
	.datac(btbframesframeblocks2tag_24),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hCCE2;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N22
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (pc_out_2 & (((\btbframes.frameblocks[1].tag [27]) # (pc_out_3)))) # (!pc_out_2 & (\btbframes.frameblocks[0].tag [27] & ((!pc_out_3))))

	.dataa(btbframesframeblocks0tag_27),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_27),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hCCE2;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N6
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (pc_out_3 & ((\btbframes.frameblocks[2].tag [26]) # ((pc_out_2)))) # (!pc_out_3 & (((!pc_out_2 & \btbframes.frameblocks[0].tag [26]))))

	.dataa(pc_out_3),
	.datab(btbframesframeblocks2tag_26),
	.datac(pc_out_2),
	.datad(btbframesframeblocks0tag_26),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hADA8;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N8
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (pc_out_2 & ((\Mux2~0_combout  & ((\btbframes.frameblocks[3].tag [26]))) # (!\Mux2~0_combout  & (\btbframes.frameblocks[1].tag [26])))) # (!pc_out_2 & (((\Mux2~0_combout ))))

	.dataa(pc_out_2),
	.datab(btbframesframeblocks1tag_26),
	.datac(btbframesframeblocks3tag_26),
	.datad(\Mux2~0_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hF588;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N6
cycloneive_lcell_comb \predicted~18 (
// Equation(s):
// predicted = (\predicted~17_combout  & (\predicted~14_combout  & (\predicted~9_combout  & \predicted~4_combout )))

	.dataa(\predicted~17_combout ),
	.datab(\predicted~14_combout ),
	.datac(\predicted~9_combout ),
	.datad(\predicted~4_combout ),
	.cin(gnd),
	.combout(predicted),
	.cout());
// synopsys translate_off
defparam \predicted~18 .lut_mask = 16'h8000;
defparam \predicted~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N18
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (pc_out_2 & (((pc_out_3)))) # (!pc_out_2 & ((pc_out_3 & (\btbframes.frameblocks[2].curr_state [1])) # (!pc_out_3 & ((\btbframes.frameblocks[0].curr_state [1])))))

	.dataa(btbframesframeblocks2curr_state_1),
	.datab(pc_out_2),
	.datac(pc_out_3),
	.datad(btbframesframeblocks0curr_state_1),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hE3E0;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N12
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (pc_out_2 & ((\Mux61~0_combout  & (\btbframes.frameblocks[3].curr_state [1])) # (!\Mux61~0_combout  & ((\btbframes.frameblocks[1].curr_state [1]))))) # (!pc_out_2 & (((\Mux61~0_combout ))))

	.dataa(btbframesframeblocks3curr_state_1),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1curr_state_1),
	.datad(\Mux61~0_combout ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hBBC0;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N8
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (pc_out_2 & (((pc_out_3) # (\btbframes.frameblocks[1].valid~q )))) # (!pc_out_2 & (\btbframes.frameblocks[0].valid~q  & (!pc_out_3)))

	.dataa(btbframesframeblocks0valid),
	.datab(pc_out_2),
	.datac(pc_out_3),
	.datad(btbframesframeblocks1valid),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hCEC2;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N4
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (\Mux0~0_combout  & ((\btbframes.frameblocks[3].valid~q ) # ((!pc_out_3)))) # (!\Mux0~0_combout  & (((pc_out_3 & \btbframes.frameblocks[2].valid~q ))))

	.dataa(btbframesframeblocks3valid),
	.datab(\Mux0~0_combout ),
	.datac(pc_out_3),
	.datad(btbframesframeblocks2valid),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hBC8C;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N8
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (\Mux4~0_combout  & (((\btbframes.frameblocks[3].tag [24])) # (!pc_out_2))) # (!\Mux4~0_combout  & (pc_out_2 & (\btbframes.frameblocks[1].tag [24])))

	.dataa(\Mux4~0_combout ),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_24),
	.datad(btbframesframeblocks3tag_24),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hEA62;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N28
cycloneive_lcell_comb \predicted~15 (
// Equation(s):
// \predicted~15_combout  = (\Mux3~1_combout  & (pc_out_29 & (\Mux4~1_combout  $ (!pc_out_28)))) # (!\Mux3~1_combout  & (!pc_out_29 & (\Mux4~1_combout  $ (!pc_out_28))))

	.dataa(\Mux3~1_combout ),
	.datab(\Mux4~1_combout ),
	.datac(pc_out_29),
	.datad(pc_out_28),
	.cin(gnd),
	.combout(\predicted~15_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~15 .lut_mask = 16'h8421;
defparam \predicted~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N10
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (\Mux1~0_combout  & ((\btbframes.frameblocks[3].tag [27]) # ((!pc_out_3)))) # (!\Mux1~0_combout  & (((\btbframes.frameblocks[2].tag [27] & pc_out_3))))

	.dataa(\Mux1~0_combout ),
	.datab(btbframesframeblocks3tag_27),
	.datac(btbframesframeblocks2tag_27),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hD8AA;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N24
cycloneive_lcell_comb \predicted~16 (
// Equation(s):
// \predicted~16_combout  = (\Mux2~1_combout  & (pc_out_30 & (\Mux1~1_combout  $ (!pc_out_31)))) # (!\Mux2~1_combout  & (!pc_out_30 & (\Mux1~1_combout  $ (!pc_out_31))))

	.dataa(\Mux2~1_combout ),
	.datab(\Mux1~1_combout ),
	.datac(pc_out_31),
	.datad(pc_out_30),
	.cin(gnd),
	.combout(\predicted~16_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~16 .lut_mask = 16'h8241;
defparam \predicted~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N30
cycloneive_lcell_comb \predicted~17 (
// Equation(s):
// \predicted~17_combout  = (!\Mux61~1_combout  & (\Mux0~1_combout  & (\predicted~15_combout  & \predicted~16_combout )))

	.dataa(\Mux61~1_combout ),
	.datab(\Mux0~1_combout ),
	.datac(\predicted~15_combout ),
	.datad(\predicted~16_combout ),
	.cin(gnd),
	.combout(\predicted~17_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~17 .lut_mask = 16'h4000;
defparam \predicted~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N20
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (pc_out_2 & ((\btbframes.frameblocks[1].tag [19]) # ((pc_out_3)))) # (!pc_out_2 & (((\btbframes.frameblocks[0].tag [19] & !pc_out_3))))

	.dataa(pc_out_2),
	.datab(btbframesframeblocks1tag_19),
	.datac(btbframesframeblocks0tag_19),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hAAD8;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N30
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (\Mux9~0_combout  & (((\btbframes.frameblocks[3].tag [19]) # (!pc_out_3)))) # (!\Mux9~0_combout  & (\btbframes.frameblocks[2].tag [19] & ((pc_out_3))))

	.dataa(btbframesframeblocks2tag_19),
	.datab(\Mux9~0_combout ),
	.datac(btbframesframeblocks3tag_19),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hE2CC;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N12
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (pc_out_3 & (((\btbframes.frameblocks[2].tag [18]) # (pc_out_2)))) # (!pc_out_3 & (\btbframes.frameblocks[0].tag [18] & ((!pc_out_2))))

	.dataa(btbframesframeblocks0tag_18),
	.datab(pc_out_3),
	.datac(btbframesframeblocks2tag_18),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hCCE2;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N14
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (pc_out_2 & ((\Mux10~0_combout  & (\btbframes.frameblocks[3].tag [18])) # (!\Mux10~0_combout  & ((\btbframes.frameblocks[1].tag [18]))))) # (!pc_out_2 & (((\Mux10~0_combout ))))

	.dataa(btbframesframeblocks3tag_18),
	.datab(btbframesframeblocks1tag_18),
	.datac(pc_out_2),
	.datad(\Mux10~0_combout ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hAFC0;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N26
cycloneive_lcell_comb \predicted~11 (
// Equation(s):
// \predicted~11_combout  = (pc_out_22 & (\Mux10~1_combout  & (\Mux9~1_combout  $ (!pc_out_23)))) # (!pc_out_22 & (!\Mux10~1_combout  & (\Mux9~1_combout  $ (!pc_out_23))))

	.dataa(pc_out_22),
	.datab(\Mux9~1_combout ),
	.datac(\Mux10~1_combout ),
	.datad(pc_out_23),
	.cin(gnd),
	.combout(\predicted~11_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~11 .lut_mask = 16'h8421;
defparam \predicted~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N12
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (pc_out_2 & (((pc_out_3)))) # (!pc_out_2 & ((pc_out_3 & ((\btbframes.frameblocks[2].tag [22]))) # (!pc_out_3 & (\btbframes.frameblocks[0].tag [22]))))

	.dataa(pc_out_2),
	.datab(btbframesframeblocks0tag_22),
	.datac(pc_out_3),
	.datad(btbframesframeblocks2tag_22),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hF4A4;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N0
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (pc_out_2 & ((\Mux6~0_combout  & (\btbframes.frameblocks[3].tag [22])) # (!\Mux6~0_combout  & ((\btbframes.frameblocks[1].tag [22]))))) # (!pc_out_2 & (((\Mux6~0_combout ))))

	.dataa(btbframesframeblocks3tag_22),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_22),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hBBC0;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N4
cycloneive_lcell_comb \predicted~13 (
// Equation(s):
// \predicted~13_combout  = (\Mux5~1_combout  & (pc_out_27 & (pc_out_26 $ (!\Mux6~1_combout )))) # (!\Mux5~1_combout  & (!pc_out_27 & (pc_out_26 $ (!\Mux6~1_combout ))))

	.dataa(\Mux5~1_combout ),
	.datab(pc_out_26),
	.datac(\Mux6~1_combout ),
	.datad(pc_out_27),
	.cin(gnd),
	.combout(\predicted~13_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~13 .lut_mask = 16'h8241;
defparam \predicted~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N16
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (\Mux7~0_combout  & (((\btbframes.frameblocks[3].tag [21])) # (!pc_out_3))) # (!\Mux7~0_combout  & (pc_out_3 & ((\btbframes.frameblocks[2].tag [21]))))

	.dataa(\Mux7~0_combout ),
	.datab(pc_out_3),
	.datac(btbframesframeblocks3tag_21),
	.datad(btbframesframeblocks2tag_21),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hE6A2;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N10
cycloneive_lcell_comb \predicted~12 (
// Equation(s):
// \predicted~12_combout  = (\Mux8~1_combout  & (pc_out_24 & (pc_out_25 $ (!\Mux7~1_combout )))) # (!\Mux8~1_combout  & (!pc_out_24 & (pc_out_25 $ (!\Mux7~1_combout ))))

	.dataa(\Mux8~1_combout ),
	.datab(pc_out_24),
	.datac(pc_out_25),
	.datad(\Mux7~1_combout ),
	.cin(gnd),
	.combout(\predicted~12_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~12 .lut_mask = 16'h9009;
defparam \predicted~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N0
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & ((\btbframes.frameblocks[1].tag [17]))) # (!pc_out_2 & (\btbframes.frameblocks[0].tag [17]))))

	.dataa(btbframesframeblocks0tag_17),
	.datab(pc_out_3),
	.datac(btbframesframeblocks1tag_17),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hFC22;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N22
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (pc_out_3 & ((\Mux11~0_combout  & ((\btbframes.frameblocks[3].tag [17]))) # (!\Mux11~0_combout  & (\btbframes.frameblocks[2].tag [17])))) # (!pc_out_3 & (((\Mux11~0_combout ))))

	.dataa(btbframesframeblocks2tag_17),
	.datab(pc_out_3),
	.datac(btbframesframeblocks3tag_17),
	.datad(\Mux11~0_combout ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hF388;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N8
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (\Mux12~0_combout  & ((\btbframes.frameblocks[3].tag [16]) # ((!pc_out_2)))) # (!\Mux12~0_combout  & (((\btbframes.frameblocks[1].tag [16] & pc_out_2))))

	.dataa(\Mux12~0_combout ),
	.datab(btbframesframeblocks3tag_16),
	.datac(btbframesframeblocks1tag_16),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hD8AA;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N6
cycloneive_lcell_comb \predicted~10 (
// Equation(s):
// \predicted~10_combout  = (pc_out_20 & (\Mux12~1_combout  & (\Mux11~1_combout  $ (!pc_out_21)))) # (!pc_out_20 & (!\Mux12~1_combout  & (\Mux11~1_combout  $ (!pc_out_21))))

	.dataa(pc_out_20),
	.datab(\Mux11~1_combout ),
	.datac(pc_out_21),
	.datad(\Mux12~1_combout ),
	.cin(gnd),
	.combout(\predicted~10_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~10 .lut_mask = 16'h8241;
defparam \predicted~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N4
cycloneive_lcell_comb \predicted~14 (
// Equation(s):
// \predicted~14_combout  = (\predicted~11_combout  & (\predicted~13_combout  & (\predicted~12_combout  & \predicted~10_combout )))

	.dataa(\predicted~11_combout ),
	.datab(\predicted~13_combout ),
	.datac(\predicted~12_combout ),
	.datad(\predicted~10_combout ),
	.cin(gnd),
	.combout(\predicted~14_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~14 .lut_mask = 16'h8000;
defparam \predicted~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N24
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (pc_out_3 & (pc_out_2)) # (!pc_out_3 & ((pc_out_2 & ((\btbframes.frameblocks[1].tag [9]))) # (!pc_out_2 & (\btbframes.frameblocks[0].tag [9]))))

	.dataa(pc_out_3),
	.datab(pc_out_2),
	.datac(btbframesframeblocks0tag_9),
	.datad(btbframesframeblocks1tag_9),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hDC98;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N10
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (pc_out_3 & ((\Mux19~0_combout  & (\btbframes.frameblocks[3].tag [9])) # (!\Mux19~0_combout  & ((\btbframes.frameblocks[2].tag [9]))))) # (!pc_out_3 & (((\Mux19~0_combout ))))

	.dataa(pc_out_3),
	.datab(btbframesframeblocks3tag_9),
	.datac(btbframesframeblocks2tag_9),
	.datad(\Mux19~0_combout ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hDDA0;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N4
cycloneive_lcell_comb \predicted~5 (
// Equation(s):
// \predicted~5_combout  = (\Mux20~1_combout  & (pc_out_12 & (\Mux19~1_combout  $ (!pc_out_13)))) # (!\Mux20~1_combout  & (!pc_out_12 & (\Mux19~1_combout  $ (!pc_out_13))))

	.dataa(\Mux20~1_combout ),
	.datab(\Mux19~1_combout ),
	.datac(pc_out_13),
	.datad(pc_out_12),
	.cin(gnd),
	.combout(\predicted~5_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~5 .lut_mask = 16'h8241;
defparam \predicted~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N6
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (\Mux16~0_combout  & (((\btbframes.frameblocks[3].tag [12])) # (!pc_out_2))) # (!\Mux16~0_combout  & (pc_out_2 & (\btbframes.frameblocks[1].tag [12])))

	.dataa(\Mux16~0_combout ),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_12),
	.datad(btbframesframeblocks3tag_12),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hEA62;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N28
cycloneive_lcell_comb \predicted~7 (
// Equation(s):
// \predicted~7_combout  = (\Mux15~1_combout  & (pc_out_17 & (pc_out_16 $ (!\Mux16~1_combout )))) # (!\Mux15~1_combout  & (!pc_out_17 & (pc_out_16 $ (!\Mux16~1_combout ))))

	.dataa(\Mux15~1_combout ),
	.datab(pc_out_17),
	.datac(pc_out_16),
	.datad(\Mux16~1_combout ),
	.cin(gnd),
	.combout(\predicted~7_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~7 .lut_mask = 16'h9009;
defparam \predicted~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N28
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (pc_out_3 & (((pc_out_2)))) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].tag [11])) # (!pc_out_2 & ((\btbframes.frameblocks[0].tag [11])))))

	.dataa(btbframesframeblocks1tag_11),
	.datab(pc_out_3),
	.datac(btbframesframeblocks0tag_11),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hEE30;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N16
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (pc_out_3 & ((\Mux17~0_combout  & ((\btbframes.frameblocks[3].tag [11]))) # (!\Mux17~0_combout  & (\btbframes.frameblocks[2].tag [11])))) # (!pc_out_3 & (((\Mux17~0_combout ))))

	.dataa(btbframesframeblocks2tag_11),
	.datab(pc_out_3),
	.datac(btbframesframeblocks3tag_11),
	.datad(\Mux17~0_combout ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hF388;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N26
cycloneive_lcell_comb \predicted~6 (
// Equation(s):
// \predicted~6_combout  = (\Mux18~1_combout  & (pc_out_14 & (pc_out_15 $ (!\Mux17~1_combout )))) # (!\Mux18~1_combout  & (!pc_out_14 & (pc_out_15 $ (!\Mux17~1_combout ))))

	.dataa(\Mux18~1_combout ),
	.datab(pc_out_14),
	.datac(pc_out_15),
	.datad(\Mux17~1_combout ),
	.cin(gnd),
	.combout(\predicted~6_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~6 .lut_mask = 16'h9009;
defparam \predicted~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N26
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (pc_out_2 & (pc_out_3)) # (!pc_out_2 & ((pc_out_3 & (\btbframes.frameblocks[2].tag [14])) # (!pc_out_3 & ((\btbframes.frameblocks[0].tag [14])))))

	.dataa(pc_out_2),
	.datab(pc_out_3),
	.datac(btbframesframeblocks2tag_14),
	.datad(btbframesframeblocks0tag_14),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hD9C8;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N12
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (pc_out_2 & ((\Mux14~0_combout  & (\btbframes.frameblocks[3].tag [14])) # (!\Mux14~0_combout  & ((\btbframes.frameblocks[1].tag [14]))))) # (!pc_out_2 & (((\Mux14~0_combout ))))

	.dataa(btbframesframeblocks3tag_14),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_14),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hBBC0;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N24
cycloneive_lcell_comb \predicted~8 (
// Equation(s):
// \predicted~8_combout  = (\Mux13~1_combout  & (pc_out_19 & (pc_out_18 $ (!\Mux14~1_combout )))) # (!\Mux13~1_combout  & (!pc_out_19 & (pc_out_18 $ (!\Mux14~1_combout ))))

	.dataa(\Mux13~1_combout ),
	.datab(pc_out_19),
	.datac(pc_out_18),
	.datad(\Mux14~1_combout ),
	.cin(gnd),
	.combout(\predicted~8_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~8 .lut_mask = 16'h9009;
defparam \predicted~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N2
cycloneive_lcell_comb \predicted~9 (
// Equation(s):
// \predicted~9_combout  = (\predicted~5_combout  & (\predicted~7_combout  & (\predicted~6_combout  & \predicted~8_combout )))

	.dataa(\predicted~5_combout ),
	.datab(\predicted~7_combout ),
	.datac(\predicted~6_combout ),
	.datad(\predicted~8_combout ),
	.cin(gnd),
	.combout(\predicted~9_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~9 .lut_mask = 16'h8000;
defparam \predicted~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N24
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (pc_out_3 & (pc_out_2)) # (!pc_out_3 & ((pc_out_2 & (\btbframes.frameblocks[1].tag [1])) # (!pc_out_2 & ((\btbframes.frameblocks[0].tag [1])))))

	.dataa(pc_out_3),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_1),
	.datad(btbframesframeblocks0tag_1),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hD9C8;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N30
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (pc_out_3 & ((\Mux27~0_combout  & (\btbframes.frameblocks[3].tag [1])) # (!\Mux27~0_combout  & ((\btbframes.frameblocks[2].tag [1]))))) # (!pc_out_3 & (\Mux27~0_combout ))

	.dataa(pc_out_3),
	.datab(\Mux27~0_combout ),
	.datac(btbframesframeblocks3tag_1),
	.datad(btbframesframeblocks2tag_1),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hE6C4;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N0
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (pc_out_2 & (pc_out_3)) # (!pc_out_2 & ((pc_out_3 & (\btbframes.frameblocks[2].tag [0])) # (!pc_out_3 & ((\btbframes.frameblocks[0].tag [0])))))

	.dataa(pc_out_2),
	.datab(pc_out_3),
	.datac(btbframesframeblocks2tag_0),
	.datad(btbframesframeblocks0tag_0),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hD9C8;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N0
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (pc_out_2 & ((\Mux28~0_combout  & (\btbframes.frameblocks[3].tag [0])) # (!\Mux28~0_combout  & ((\btbframes.frameblocks[1].tag [0]))))) # (!pc_out_2 & (((\Mux28~0_combout ))))

	.dataa(btbframesframeblocks3tag_0),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_0),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hBBC0;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N20
cycloneive_lcell_comb \predicted~0 (
// Equation(s):
// \predicted~0_combout  = (pc_out_4 & (\Mux28~1_combout  & (pc_out_5 $ (!\Mux27~1_combout )))) # (!pc_out_4 & (!\Mux28~1_combout  & (pc_out_5 $ (!\Mux27~1_combout ))))

	.dataa(pc_out_4),
	.datab(pc_out_5),
	.datac(\Mux27~1_combout ),
	.datad(\Mux28~1_combout ),
	.cin(gnd),
	.combout(\predicted~0_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~0 .lut_mask = 16'h8241;
defparam \predicted~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N6
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (pc_out_3 & (((\btbframes.frameblocks[2].tag [4]) # (pc_out_2)))) # (!pc_out_3 & (\btbframes.frameblocks[0].tag [4] & ((!pc_out_2))))

	.dataa(pc_out_3),
	.datab(btbframesframeblocks0tag_4),
	.datac(btbframesframeblocks2tag_4),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hAAE4;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N24
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (pc_out_2 & ((\Mux24~0_combout  & ((\btbframes.frameblocks[3].tag [4]))) # (!\Mux24~0_combout  & (\btbframes.frameblocks[1].tag [4])))) # (!pc_out_2 & (((\Mux24~0_combout ))))

	.dataa(btbframesframeblocks1tag_4),
	.datab(pc_out_2),
	.datac(btbframesframeblocks3tag_4),
	.datad(\Mux24~0_combout ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hF388;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N22
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (pc_out_2 & (((pc_out_3) # (\btbframes.frameblocks[1].tag [5])))) # (!pc_out_2 & (\btbframes.frameblocks[0].tag [5] & (!pc_out_3)))

	.dataa(pc_out_2),
	.datab(btbframesframeblocks0tag_5),
	.datac(pc_out_3),
	.datad(btbframesframeblocks1tag_5),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hAEA4;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N20
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (pc_out_3 & ((\Mux23~0_combout  & (\btbframes.frameblocks[3].tag [5])) # (!\Mux23~0_combout  & ((\btbframes.frameblocks[2].tag [5]))))) # (!pc_out_3 & (((\Mux23~0_combout ))))

	.dataa(pc_out_3),
	.datab(btbframesframeblocks3tag_5),
	.datac(\Mux23~0_combout ),
	.datad(btbframesframeblocks2tag_5),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hDAD0;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N4
cycloneive_lcell_comb \predicted~2 (
// Equation(s):
// \predicted~2_combout  = (pc_out_8 & (\Mux24~1_combout  & (pc_out_9 $ (!\Mux23~1_combout )))) # (!pc_out_8 & (!\Mux24~1_combout  & (pc_out_9 $ (!\Mux23~1_combout ))))

	.dataa(pc_out_8),
	.datab(pc_out_9),
	.datac(\Mux24~1_combout ),
	.datad(\Mux23~1_combout ),
	.cin(gnd),
	.combout(\predicted~2_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~2 .lut_mask = 16'h8421;
defparam \predicted~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N16
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (pc_out_3 & (((\btbframes.frameblocks[2].tag [6]) # (pc_out_2)))) # (!pc_out_3 & (\btbframes.frameblocks[0].tag [6] & ((!pc_out_2))))

	.dataa(btbframesframeblocks0tag_6),
	.datab(btbframesframeblocks2tag_6),
	.datac(pc_out_3),
	.datad(pc_out_2),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hF0CA;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N14
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (pc_out_2 & ((\Mux22~0_combout  & (\btbframes.frameblocks[3].tag [6])) # (!\Mux22~0_combout  & ((\btbframes.frameblocks[1].tag [6]))))) # (!pc_out_2 & (((\Mux22~0_combout ))))

	.dataa(btbframesframeblocks3tag_6),
	.datab(pc_out_2),
	.datac(btbframesframeblocks1tag_6),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hBBC0;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N28
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (\Mux21~0_combout  & (((\btbframes.frameblocks[3].tag [7]) # (!pc_out_3)))) # (!\Mux21~0_combout  & (\btbframes.frameblocks[2].tag [7] & ((pc_out_3))))

	.dataa(\Mux21~0_combout ),
	.datab(btbframesframeblocks2tag_7),
	.datac(btbframesframeblocks3tag_7),
	.datad(pc_out_3),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hE4AA;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N30
cycloneive_lcell_comb \predicted~3 (
// Equation(s):
// \predicted~3_combout  = (pc_out_11 & (\Mux21~1_combout  & (pc_out_10 $ (!\Mux22~1_combout )))) # (!pc_out_11 & (!\Mux21~1_combout  & (pc_out_10 $ (!\Mux22~1_combout ))))

	.dataa(pc_out_11),
	.datab(pc_out_10),
	.datac(\Mux22~1_combout ),
	.datad(\Mux21~1_combout ),
	.cin(gnd),
	.combout(\predicted~3_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~3 .lut_mask = 16'h8241;
defparam \predicted~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N22
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (pc_out_2 & (pc_out_3)) # (!pc_out_2 & ((pc_out_3 & (\btbframes.frameblocks[2].tag [2])) # (!pc_out_3 & ((\btbframes.frameblocks[0].tag [2])))))

	.dataa(pc_out_2),
	.datab(pc_out_3),
	.datac(btbframesframeblocks2tag_2),
	.datad(btbframesframeblocks0tag_2),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hD9C8;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N2
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (pc_out_2 & ((\Mux26~0_combout  & ((\btbframes.frameblocks[3].tag [2]))) # (!\Mux26~0_combout  & (\btbframes.frameblocks[1].tag [2])))) # (!pc_out_2 & (((\Mux26~0_combout ))))

	.dataa(btbframesframeblocks1tag_2),
	.datab(btbframesframeblocks3tag_2),
	.datac(pc_out_2),
	.datad(\Mux26~0_combout ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hCFA0;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N6
cycloneive_lcell_comb \predicted~1 (
// Equation(s):
// \predicted~1_combout  = (\Mux25~1_combout  & (pc_out_7 & (pc_out_6 $ (!\Mux26~1_combout )))) # (!\Mux25~1_combout  & (!pc_out_7 & (pc_out_6 $ (!\Mux26~1_combout ))))

	.dataa(\Mux25~1_combout ),
	.datab(pc_out_6),
	.datac(\Mux26~1_combout ),
	.datad(pc_out_7),
	.cin(gnd),
	.combout(\predicted~1_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~1 .lut_mask = 16'h8241;
defparam \predicted~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N24
cycloneive_lcell_comb \predicted~4 (
// Equation(s):
// \predicted~4_combout  = (\predicted~0_combout  & (\predicted~2_combout  & (\predicted~3_combout  & \predicted~1_combout )))

	.dataa(\predicted~0_combout ),
	.datab(\predicted~2_combout ),
	.datac(\predicted~3_combout ),
	.datad(\predicted~1_combout ),
	.cin(gnd),
	.combout(\predicted~4_combout ),
	.cout());
// synopsys translate_off
defparam \predicted~4 .lut_mask = 16'h8000;
defparam \predicted~4 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module control_unit (
	instruction_D_31,
	instruction_D_28,
	instruction_D_30,
	instruction_D_29,
	instruction_D_27,
	instruction_D_26,
	Decoder1,
	Decoder11,
	Equal3,
	Equal31,
	instruction_D_5,
	instruction_D_0,
	instruction_D_3,
	instruction_D_2,
	instruction_D_1,
	WideOr2,
	instruction_D_4,
	WideOr7,
	WideOr6,
	WideOr1,
	WideOr5,
	WideOr8,
	WideOr4,
	Decoder0,
	devpor,
	devclrn,
	devoe);
input 	instruction_D_31;
input 	instruction_D_28;
input 	instruction_D_30;
input 	instruction_D_29;
input 	instruction_D_27;
input 	instruction_D_26;
output 	Decoder1;
output 	Decoder11;
output 	Equal3;
output 	Equal31;
input 	instruction_D_5;
input 	instruction_D_0;
input 	instruction_D_3;
input 	instruction_D_2;
input 	instruction_D_1;
output 	WideOr2;
input 	instruction_D_4;
output 	WideOr7;
output 	WideOr6;
output 	WideOr1;
output 	WideOr5;
output 	WideOr8;
output 	WideOr4;
output 	Decoder0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Equal3~0_combout ;
wire \Decoder0~0_combout ;


// Location: LCCOMB_X63_Y38_N10
cycloneive_lcell_comb \Decoder1~0 (
// Equation(s):
// Decoder1 = (instruction_D[26] & (instruction_D[29] & instruction_D[27]))

	.dataa(instruction_D_26),
	.datab(gnd),
	.datac(instruction_D_29),
	.datad(instruction_D_27),
	.cin(gnd),
	.combout(Decoder1),
	.cout());
// synopsys translate_off
defparam \Decoder1~0 .lut_mask = 16'hA000;
defparam \Decoder1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N0
cycloneive_lcell_comb \Decoder1~1 (
// Equation(s):
// Decoder11 = (instruction_D[31] & (instruction_D[30] & (instruction_D[28] & Decoder1)))

	.dataa(instruction_D_31),
	.datab(instruction_D_30),
	.datac(instruction_D_28),
	.datad(Decoder1),
	.cin(gnd),
	.combout(Decoder11),
	.cout());
// synopsys translate_off
defparam \Decoder1~1 .lut_mask = 16'h8000;
defparam \Decoder1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N2
cycloneive_lcell_comb \Equal3~1 (
// Equation(s):
// Equal3 = (!instruction_D[29] & !instruction_D[28])

	.dataa(gnd),
	.datab(instruction_D_29),
	.datac(instruction_D_28),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal3),
	.cout());
// synopsys translate_off
defparam \Equal3~1 .lut_mask = 16'h0303;
defparam \Equal3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N2
cycloneive_lcell_comb \Equal3~2 (
// Equation(s):
// Equal31 = (!instruction_D[26] & (!instruction_D[27] & (\Equal3~0_combout  & Equal3)))

	.dataa(instruction_D_26),
	.datab(instruction_D_27),
	.datac(\Equal3~0_combout ),
	.datad(Equal3),
	.cin(gnd),
	.combout(Equal31),
	.cout());
// synopsys translate_off
defparam \Equal3~2 .lut_mask = 16'h1000;
defparam \Equal3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N20
cycloneive_lcell_comb \WideOr2~0 (
// Equation(s):
// WideOr2 = (instruction_D[2] & (!instruction_D[3] & ((instruction_D[0])))) # (!instruction_D[2] & (instruction_D[1] & ((instruction_D[0]) # (!instruction_D[3]))))

	.dataa(instruction_D_2),
	.datab(instruction_D_3),
	.datac(instruction_D_1),
	.datad(instruction_D_0),
	.cin(gnd),
	.combout(WideOr2),
	.cout());
// synopsys translate_off
defparam \WideOr2~0 .lut_mask = 16'h7210;
defparam \WideOr2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N4
cycloneive_lcell_comb \WideOr7~0 (
// Equation(s):
// WideOr7 = (instruction_D[29] & (instruction_D[26] & (instruction_D[28] $ (instruction_D[27])))) # (!instruction_D[29] & (((instruction_D[28] & !instruction_D[27]))))

	.dataa(instruction_D_26),
	.datab(instruction_D_29),
	.datac(instruction_D_28),
	.datad(instruction_D_27),
	.cin(gnd),
	.combout(WideOr7),
	.cout());
// synopsys translate_off
defparam \WideOr7~0 .lut_mask = 16'h08B0;
defparam \WideOr7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N0
cycloneive_lcell_comb \WideOr6~0 (
// Equation(s):
// WideOr6 = (instruction_D[28] & ((instruction_D[27] & (instruction_D[29] & !instruction_D[26])) # (!instruction_D[27] & (!instruction_D[29])))) # (!instruction_D[28] & (((instruction_D[29]))))

	.dataa(instruction_D_28),
	.datab(instruction_D_27),
	.datac(instruction_D_29),
	.datad(instruction_D_26),
	.cin(gnd),
	.combout(WideOr6),
	.cout());
// synopsys translate_off
defparam \WideOr6~0 .lut_mask = 16'h52D2;
defparam \WideOr6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N0
cycloneive_lcell_comb \WideOr1~0 (
// Equation(s):
// WideOr1 = (instruction_D[4]) # ((instruction_D[2] & ((instruction_D[3]) # (!instruction_D[1]))) # (!instruction_D[2] & (instruction_D[3] & !instruction_D[1])))

	.dataa(instruction_D_2),
	.datab(instruction_D_3),
	.datac(instruction_D_1),
	.datad(instruction_D_4),
	.cin(gnd),
	.combout(WideOr1),
	.cout());
// synopsys translate_off
defparam \WideOr1~0 .lut_mask = 16'hFF8E;
defparam \WideOr1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N30
cycloneive_lcell_comb \WideOr5~0 (
// Equation(s):
// WideOr5 = (instruction_D[28] & (instruction_D[29] & ((!instruction_D[26]) # (!instruction_D[27]))))

	.dataa(instruction_D_28),
	.datab(instruction_D_27),
	.datac(instruction_D_29),
	.datad(instruction_D_26),
	.cin(gnd),
	.combout(WideOr5),
	.cout());
// synopsys translate_off
defparam \WideOr5~0 .lut_mask = 16'h20A0;
defparam \WideOr5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N18
cycloneive_lcell_comb \WideOr8~0 (
// Equation(s):
// WideOr8 = (instruction_D[31] & (instruction_D[26] & (instruction_D[27]))) # (!instruction_D[31] & (((instruction_D[29]))))

	.dataa(instruction_D_26),
	.datab(instruction_D_27),
	.datac(instruction_D_29),
	.datad(instruction_D_31),
	.cin(gnd),
	.combout(WideOr8),
	.cout());
// synopsys translate_off
defparam \WideOr8~0 .lut_mask = 16'h88F0;
defparam \WideOr8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N22
cycloneive_lcell_comb \WideOr4~0 (
// Equation(s):
// WideOr4 = (instruction_D[31] & (((instruction_D[28]) # (!instruction_D[27])) # (!instruction_D[26])))

	.dataa(instruction_D_26),
	.datab(instruction_D_27),
	.datac(instruction_D_31),
	.datad(instruction_D_28),
	.cin(gnd),
	.combout(WideOr4),
	.cout());
// synopsys translate_off
defparam \WideOr4~0 .lut_mask = 16'hF070;
defparam \WideOr4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N8
cycloneive_lcell_comb \Decoder0~1 (
// Equation(s):
// Decoder0 = (instruction_D[1]) # ((\Decoder0~0_combout ) # (!instruction_D[3]))

	.dataa(instruction_D_1),
	.datab(instruction_D_3),
	.datac(gnd),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(Decoder0),
	.cout());
// synopsys translate_off
defparam \Decoder0~1 .lut_mask = 16'hFFBB;
defparam \Decoder0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N4
cycloneive_lcell_comb \Equal3~0 (
// Equation(s):
// \Equal3~0_combout  = (!instruction_D[30] & !instruction_D[31])

	.dataa(gnd),
	.datab(instruction_D_30),
	.datac(gnd),
	.datad(instruction_D_31),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~0 .lut_mask = 16'h0033;
defparam \Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N10
cycloneive_lcell_comb \Decoder0~0 (
// Equation(s):
// \Decoder0~0_combout  = (instruction_D[2]) # ((instruction_D[0]) # ((instruction_D[4]) # (instruction_D[5])))

	.dataa(instruction_D_2),
	.datab(instruction_D_0),
	.datac(instruction_D_4),
	.datad(instruction_D_5),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~0 .lut_mask = 16'hFFFE;
defparam \Decoder0~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module forwarding_unit (
	dREN_M,
	Equal4,
	op_EX_1,
	op_EX_0,
	Equal41,
	instruction_EX_16,
	instruction_EX_17,
	wsel_M_1,
	wsel_M_0,
	instruction_EX_18,
	instruction_EX_19,
	wsel_M_3,
	wsel_M_2,
	instruction_EX_20,
	wsel_M_4,
	Equal0,
	instruction_EX_22,
	instruction_EX_21,
	instruction_EX_24,
	instruction_EX_23,
	instruction_EX_25,
	fuifforward_A_0,
	wsel_WB_1,
	wsel_WB_0,
	wsel_WB_3,
	wsel_WB_2,
	wsel_WB_4,
	fuifforward_A_1,
	fuifbubble_lw_f,
	regWrite_M,
	forward_B,
	beq_EX,
	bne_EX,
	forward_B1,
	Equal5,
	regWrite_WB,
	fuifforward_B_1,
	fuifforward_B_11,
	Equal3,
	fuifforward_A_01,
	Equal31,
	fuifforward_A_11,
	devpor,
	devclrn,
	devoe);
input 	dREN_M;
input 	Equal4;
input 	op_EX_1;
input 	op_EX_0;
input 	Equal41;
input 	instruction_EX_16;
input 	instruction_EX_17;
input 	wsel_M_1;
input 	wsel_M_0;
input 	instruction_EX_18;
input 	instruction_EX_19;
input 	wsel_M_3;
input 	wsel_M_2;
input 	instruction_EX_20;
input 	wsel_M_4;
output 	Equal0;
input 	instruction_EX_22;
input 	instruction_EX_21;
input 	instruction_EX_24;
input 	instruction_EX_23;
input 	instruction_EX_25;
output 	fuifforward_A_0;
input 	wsel_WB_1;
input 	wsel_WB_0;
input 	wsel_WB_3;
input 	wsel_WB_2;
input 	wsel_WB_4;
output 	fuifforward_A_1;
output 	fuifbubble_lw_f;
input 	regWrite_M;
output 	forward_B;
input 	beq_EX;
input 	bne_EX;
output 	forward_B1;
output 	Equal5;
input 	regWrite_WB;
output 	fuifforward_B_1;
output 	fuifforward_B_11;
output 	Equal3;
output 	fuifforward_A_01;
output 	Equal31;
output 	fuifforward_A_11;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \fuif.forward_A[0]~0_combout ;
wire \fuif.forward_A[0]~1_combout ;
wire \fuif.forward_A[1]~3_combout ;
wire \fuif.forward_A[1]~4_combout ;
wire \fuif.bubble_lw_f~3_combout ;
wire \Equal0~3_combout ;
wire \Equal5~0_combout ;
wire \fuif.forward_B[1]~1_combout ;
wire \fuif.forward_B[1]~2_combout ;
wire \forward_B~2_combout ;
wire \fuif.forward_B[1]~0_combout ;


// Location: LCCOMB_X62_Y35_N24
cycloneive_lcell_comb \Equal0~2 (
// Equation(s):
// Equal0 = (\Equal0~0_combout  & (\Equal0~1_combout  & (wsel_M[4] $ (!instruction_EX[20]))))

	.dataa(\Equal0~0_combout ),
	.datab(wsel_M_4),
	.datac(instruction_EX_20),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~2 .lut_mask = 16'h8200;
defparam \Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N2
cycloneive_lcell_comb \fuif.forward_A[0]~2 (
// Equation(s):
// fuifforward_A_0 = (\fuif.forward_A[0]~0_combout  & (\fuif.forward_A[0]~1_combout  & (instruction_EX[25] $ (!wsel_M[4]))))

	.dataa(instruction_EX_25),
	.datab(wsel_M_4),
	.datac(\fuif.forward_A[0]~0_combout ),
	.datad(\fuif.forward_A[0]~1_combout ),
	.cin(gnd),
	.combout(fuifforward_A_0),
	.cout());
// synopsys translate_off
defparam \fuif.forward_A[0]~2 .lut_mask = 16'h9000;
defparam \fuif.forward_A[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N26
cycloneive_lcell_comb \fuif.forward_A[1]~5 (
// Equation(s):
// fuifforward_A_1 = (\fuif.forward_A[1]~3_combout  & (\fuif.forward_A[1]~4_combout  & (instruction_EX[25] $ (!wsel_WB[4]))))

	.dataa(instruction_EX_25),
	.datab(wsel_WB_4),
	.datac(\fuif.forward_A[1]~3_combout ),
	.datad(\fuif.forward_A[1]~4_combout ),
	.cin(gnd),
	.combout(fuifforward_A_1),
	.cout());
// synopsys translate_off
defparam \fuif.forward_A[1]~5 .lut_mask = 16'h9000;
defparam \fuif.forward_A[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N20
cycloneive_lcell_comb \fuif.bubble_lw_f~2 (
// Equation(s):
// fuifbubble_lw_f = (dREN_M1 & ((fuifforward_A_0) # ((fuifforward_A_1) # (\fuif.bubble_lw_f~3_combout ))))

	.dataa(dREN_M),
	.datab(fuifforward_A_0),
	.datac(fuifforward_A_1),
	.datad(\fuif.bubble_lw_f~3_combout ),
	.cin(gnd),
	.combout(fuifbubble_lw_f),
	.cout());
// synopsys translate_off
defparam \fuif.bubble_lw_f~2 .lut_mask = 16'hAAA8;
defparam \fuif.bubble_lw_f~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N14
cycloneive_lcell_comb \forward_B~0 (
// Equation(s):
// forward_B = (\regWrite_M~q  & (!\Equal0~3_combout  & (\Equal0~0_combout  & \Equal0~1_combout )))

	.dataa(regWrite_M),
	.datab(\Equal0~3_combout ),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(forward_B),
	.cout());
// synopsys translate_off
defparam \forward_B~0 .lut_mask = 16'h2000;
defparam \forward_B~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N12
cycloneive_lcell_comb \forward_B~1 (
// Equation(s):
// forward_B1 = (!\bne_EX~q  & (!\beq_EX~q  & ((!\Equal4~1_combout ) # (!\Equal4~0_combout ))))

	.dataa(Equal4),
	.datab(bne_EX),
	.datac(Equal41),
	.datad(beq_EX),
	.cin(gnd),
	.combout(forward_B1),
	.cout());
// synopsys translate_off
defparam \forward_B~1 .lut_mask = 16'h0013;
defparam \forward_B~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N18
cycloneive_lcell_comb \Equal5~1 (
// Equation(s):
// Equal5 = (!instruction_EX[20] & (!instruction_EX[19] & (!instruction_EX[16] & \Equal5~0_combout )))

	.dataa(instruction_EX_20),
	.datab(instruction_EX_19),
	.datac(instruction_EX_16),
	.datad(\Equal5~0_combout ),
	.cin(gnd),
	.combout(Equal5),
	.cout());
// synopsys translate_off
defparam \Equal5~1 .lut_mask = 16'h0100;
defparam \Equal5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N2
cycloneive_lcell_comb \fuif.forward_B[1]~3 (
// Equation(s):
// fuifforward_B_1 = (\fuif.forward_B[1]~1_combout  & (\fuif.forward_B[1]~2_combout  & (instruction_EX[20] $ (!wsel_WB[4]))))

	.dataa(instruction_EX_20),
	.datab(\fuif.forward_B[1]~1_combout ),
	.datac(wsel_WB_4),
	.datad(\fuif.forward_B[1]~2_combout ),
	.cin(gnd),
	.combout(fuifforward_B_1),
	.cout());
// synopsys translate_off
defparam \fuif.forward_B[1]~3 .lut_mask = 16'h8400;
defparam \fuif.forward_B[1]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N28
cycloneive_lcell_comb \fuif.forward_B[1]~4 (
// Equation(s):
// fuifforward_B_11 = (\fuif.forward_B[1]~0_combout  & (!Equal5 & (!forward_B & fuifforward_B_1)))

	.dataa(\fuif.forward_B[1]~0_combout ),
	.datab(Equal5),
	.datac(forward_B),
	.datad(fuifforward_B_1),
	.cin(gnd),
	.combout(fuifforward_B_11),
	.cout());
// synopsys translate_off
defparam \fuif.forward_B[1]~4 .lut_mask = 16'h0200;
defparam \fuif.forward_B[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N26
cycloneive_lcell_comb \Equal3~0 (
// Equation(s):
// Equal3 = (!instruction_EX[22] & (!instruction_EX[23] & (!instruction_EX[25] & !instruction_EX[24])))

	.dataa(instruction_EX_22),
	.datab(instruction_EX_23),
	.datac(instruction_EX_25),
	.datad(instruction_EX_24),
	.cin(gnd),
	.combout(Equal3),
	.cout());
// synopsys translate_off
defparam \Equal3~0 .lut_mask = 16'h0001;
defparam \Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N4
cycloneive_lcell_comb \fuif.forward_A[0]~6 (
// Equation(s):
// fuifforward_A_01 = (\regWrite_M~q  & (fuifforward_A_0 & ((instruction_EX[21]) # (!Equal3))))

	.dataa(regWrite_M),
	.datab(instruction_EX_21),
	.datac(Equal3),
	.datad(fuifforward_A_0),
	.cin(gnd),
	.combout(fuifforward_A_01),
	.cout());
// synopsys translate_off
defparam \fuif.forward_A[0]~6 .lut_mask = 16'h8A00;
defparam \fuif.forward_A[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N6
cycloneive_lcell_comb \Equal3~1 (
// Equation(s):
// Equal31 = (!instruction_EX[21] & Equal3)

	.dataa(gnd),
	.datab(instruction_EX_21),
	.datac(Equal3),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal31),
	.cout());
// synopsys translate_off
defparam \Equal3~1 .lut_mask = 16'h3030;
defparam \Equal3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N16
cycloneive_lcell_comb \fuif.forward_A[1]~7 (
// Equation(s):
// fuifforward_A_11 = (fuifforward_A_1 & (\regWrite_WB~q  & (!fuifforward_A_01 & !Equal31)))

	.dataa(fuifforward_A_1),
	.datab(regWrite_WB),
	.datac(fuifforward_A_01),
	.datad(Equal31),
	.cin(gnd),
	.combout(fuifforward_A_11),
	.cout());
// synopsys translate_off
defparam \fuif.forward_A[1]~7 .lut_mask = 16'h0008;
defparam \fuif.forward_A[1]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N0
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (instruction_EX[17] & (wsel_M[1] & (wsel_M[0] $ (!instruction_EX[16])))) # (!instruction_EX[17] & (!wsel_M[1] & (wsel_M[0] $ (!instruction_EX[16]))))

	.dataa(instruction_EX_17),
	.datab(wsel_M_0),
	.datac(wsel_M_1),
	.datad(instruction_EX_16),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h8421;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N10
cycloneive_lcell_comb \Equal0~1 (
// Equation(s):
// \Equal0~1_combout  = (wsel_M[3] & (instruction_EX[19] & (instruction_EX[18] $ (!wsel_M[2])))) # (!wsel_M[3] & (!instruction_EX[19] & (instruction_EX[18] $ (!wsel_M[2]))))

	.dataa(wsel_M_3),
	.datab(instruction_EX_18),
	.datac(wsel_M_2),
	.datad(instruction_EX_19),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~1 .lut_mask = 16'h8241;
defparam \Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N30
cycloneive_lcell_comb \fuif.forward_A[0]~0 (
// Equation(s):
// \fuif.forward_A[0]~0_combout  = (wsel_M[0] & (instruction_EX[21] & (wsel_M[1] $ (!instruction_EX[22])))) # (!wsel_M[0] & (!instruction_EX[21] & (wsel_M[1] $ (!instruction_EX[22]))))

	.dataa(wsel_M_0),
	.datab(instruction_EX_21),
	.datac(wsel_M_1),
	.datad(instruction_EX_22),
	.cin(gnd),
	.combout(\fuif.forward_A[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \fuif.forward_A[0]~0 .lut_mask = 16'h9009;
defparam \fuif.forward_A[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N24
cycloneive_lcell_comb \fuif.forward_A[0]~1 (
// Equation(s):
// \fuif.forward_A[0]~1_combout  = (wsel_M[2] & (instruction_EX[23] & (wsel_M[3] $ (!instruction_EX[24])))) # (!wsel_M[2] & (!instruction_EX[23] & (wsel_M[3] $ (!instruction_EX[24]))))

	.dataa(wsel_M_2),
	.datab(wsel_M_3),
	.datac(instruction_EX_24),
	.datad(instruction_EX_23),
	.cin(gnd),
	.combout(\fuif.forward_A[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \fuif.forward_A[0]~1 .lut_mask = 16'h8241;
defparam \fuif.forward_A[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N0
cycloneive_lcell_comb \fuif.forward_A[1]~3 (
// Equation(s):
// \fuif.forward_A[1]~3_combout  = (wsel_WB[0] & (instruction_EX[21] & (instruction_EX[22] $ (!wsel_WB[1])))) # (!wsel_WB[0] & (!instruction_EX[21] & (instruction_EX[22] $ (!wsel_WB[1]))))

	.dataa(wsel_WB_0),
	.datab(instruction_EX_22),
	.datac(wsel_WB_1),
	.datad(instruction_EX_21),
	.cin(gnd),
	.combout(\fuif.forward_A[1]~3_combout ),
	.cout());
// synopsys translate_off
defparam \fuif.forward_A[1]~3 .lut_mask = 16'h8241;
defparam \fuif.forward_A[1]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N20
cycloneive_lcell_comb \fuif.forward_A[1]~4 (
// Equation(s):
// \fuif.forward_A[1]~4_combout  = (wsel_WB[3] & (instruction_EX[24] & (wsel_WB[2] $ (!instruction_EX[23])))) # (!wsel_WB[3] & (!instruction_EX[24] & (wsel_WB[2] $ (!instruction_EX[23]))))

	.dataa(wsel_WB_3),
	.datab(wsel_WB_2),
	.datac(instruction_EX_24),
	.datad(instruction_EX_23),
	.cin(gnd),
	.combout(\fuif.forward_A[1]~4_combout ),
	.cout());
// synopsys translate_off
defparam \fuif.forward_A[1]~4 .lut_mask = 16'h8421;
defparam \fuif.forward_A[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N18
cycloneive_lcell_comb \fuif.bubble_lw_f~3 (
// Equation(s):
// \fuif.bubble_lw_f~3_combout  = (\Equal4~0_combout  & (Equal0 & (op_EX[1] & op_EX[0])))

	.dataa(Equal4),
	.datab(Equal0),
	.datac(op_EX_1),
	.datad(op_EX_0),
	.cin(gnd),
	.combout(\fuif.bubble_lw_f~3_combout ),
	.cout());
// synopsys translate_off
defparam \fuif.bubble_lw_f~3 .lut_mask = 16'h8000;
defparam \fuif.bubble_lw_f~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N0
cycloneive_lcell_comb \Equal0~3 (
// Equation(s):
// \Equal0~3_combout  = instruction_EX[20] $ (wsel_M[4])

	.dataa(gnd),
	.datab(instruction_EX_20),
	.datac(gnd),
	.datad(wsel_M_4),
	.cin(gnd),
	.combout(\Equal0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~3 .lut_mask = 16'h33CC;
defparam \Equal0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N12
cycloneive_lcell_comb \Equal5~0 (
// Equation(s):
// \Equal5~0_combout  = (!instruction_EX[18] & !instruction_EX[17])

	.dataa(gnd),
	.datab(gnd),
	.datac(instruction_EX_18),
	.datad(instruction_EX_17),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal5~0 .lut_mask = 16'h000F;
defparam \Equal5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N8
cycloneive_lcell_comb \fuif.forward_B[1]~1 (
// Equation(s):
// \fuif.forward_B[1]~1_combout  = (wsel_WB[0] & (instruction_EX[16] & (wsel_WB[1] $ (!instruction_EX[17])))) # (!wsel_WB[0] & (!instruction_EX[16] & (wsel_WB[1] $ (!instruction_EX[17]))))

	.dataa(wsel_WB_0),
	.datab(wsel_WB_1),
	.datac(instruction_EX_17),
	.datad(instruction_EX_16),
	.cin(gnd),
	.combout(\fuif.forward_B[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \fuif.forward_B[1]~1 .lut_mask = 16'h8241;
defparam \fuif.forward_B[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N18
cycloneive_lcell_comb \fuif.forward_B[1]~2 (
// Equation(s):
// \fuif.forward_B[1]~2_combout  = (wsel_WB[3] & (instruction_EX[19] & (wsel_WB[2] $ (!instruction_EX[18])))) # (!wsel_WB[3] & (!instruction_EX[19] & (wsel_WB[2] $ (!instruction_EX[18]))))

	.dataa(wsel_WB_3),
	.datab(wsel_WB_2),
	.datac(instruction_EX_18),
	.datad(instruction_EX_19),
	.cin(gnd),
	.combout(\fuif.forward_B[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \fuif.forward_B[1]~2 .lut_mask = 16'h8241;
defparam \fuif.forward_B[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N16
cycloneive_lcell_comb \forward_B~2 (
// Equation(s):
// \forward_B~2_combout  = (!\bne_EX~q  & !\beq_EX~q )

	.dataa(gnd),
	.datab(gnd),
	.datac(bne_EX),
	.datad(beq_EX),
	.cin(gnd),
	.combout(\forward_B~2_combout ),
	.cout());
// synopsys translate_off
defparam \forward_B~2 .lut_mask = 16'h000F;
defparam \forward_B~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N22
cycloneive_lcell_comb \fuif.forward_B[1]~0 (
// Equation(s):
// \fuif.forward_B[1]~0_combout  = (\regWrite_WB~q  & (((\Equal4~0_combout  & \Equal4~1_combout )) # (!\forward_B~2_combout )))

	.dataa(Equal4),
	.datab(regWrite_WB),
	.datac(Equal41),
	.datad(\forward_B~2_combout ),
	.cin(gnd),
	.combout(\fuif.forward_B[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \fuif.forward_B[1]~0 .lut_mask = 16'h80CC;
defparam \fuif.forward_B[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module program_counter (
	pc_out_3,
	pc_out_2,
	pc_out_5,
	pc_out_4,
	pc_out_7,
	pc_out_6,
	pc_out_9,
	pc_out_8,
	pc_out_11,
	pc_out_10,
	pc_out_13,
	pc_out_12,
	pc_out_15,
	pc_out_14,
	pc_out_17,
	pc_out_16,
	pc_out_19,
	pc_out_18,
	pc_out_21,
	pc_out_20,
	pc_out_23,
	pc_out_22,
	pc_out_25,
	pc_out_24,
	pc_out_27,
	pc_out_26,
	predicted_M,
	pc_plus_4_2,
	pc_plus_4_3,
	pc_plus_4_4,
	pc_plus_4_5,
	pc_plus_4_6,
	pc_plus_4_7,
	pc_plus_4_8,
	pc_plus_4_9,
	pc_plus_4_10,
	pc_plus_4_11,
	pc_plus_4_12,
	pc_plus_4_13,
	pc_plus_4_14,
	pc_plus_4_15,
	pc_plus_4_16,
	pc_plus_4_17,
	pc_plus_4_18,
	pc_plus_4_19,
	pc_plus_4_20,
	pc_plus_4_21,
	pc_plus_4_22,
	pc_plus_4_23,
	pc_plus_4_24,
	pc_plus_4_25,
	pc_plus_4_26,
	pc_plus_4_27,
	pc_out_1,
	pc_out_0,
	pc_out_29,
	pc_out_28,
	pc_out_31,
	pc_out_30,
	j_M,
	jal_M,
	branch_or_jump,
	branch_taken,
	jr_M,
	branch_or_jump1,
	predicted,
	pc_next,
	pc_next_1,
	pc_next_0,
	pc_next_3,
	pc_next_31,
	comb,
	pc_next_2,
	pc_next_21,
	pc_next_5,
	pc_next_51,
	pc_next_4,
	pc_next_41,
	pc_next_7,
	pc_next_71,
	pc_next_6,
	pc_next_61,
	pc_next_9,
	pc_next_91,
	pc_next_8,
	pc_next_81,
	pc_next_11,
	pc_next_111,
	pc_next_10,
	pc_next_101,
	pc_next_13,
	pc_next_131,
	pc_next_12,
	pc_next_121,
	pc_next_15,
	pc_next_151,
	pc_next_14,
	pc_next_141,
	pc_next_17,
	pc_next_171,
	pc_next_16,
	pc_next_161,
	pc_next_19,
	pc_next_191,
	pc_next_18,
	pc_next_181,
	pc_next_211,
	pc_next_212,
	pc_next_20,
	pc_next_201,
	pc_next_23,
	pc_next_231,
	pc_next_22,
	pc_next_221,
	pc_next_25,
	pc_next_251,
	pc_next_24,
	pc_next_241,
	pc_next_27,
	pc_next_271,
	pc_next_26,
	pc_next_261,
	pc_out_291,
	pc_out_292,
	pc_next_29,
	pc_next_28,
	pc_next_311,
	pc_next_30,
	comb1,
	pc_out_101,
	nRST,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	pc_out_3;
output 	pc_out_2;
output 	pc_out_5;
output 	pc_out_4;
output 	pc_out_7;
output 	pc_out_6;
output 	pc_out_9;
output 	pc_out_8;
output 	pc_out_11;
output 	pc_out_10;
output 	pc_out_13;
output 	pc_out_12;
output 	pc_out_15;
output 	pc_out_14;
output 	pc_out_17;
output 	pc_out_16;
output 	pc_out_19;
output 	pc_out_18;
output 	pc_out_21;
output 	pc_out_20;
output 	pc_out_23;
output 	pc_out_22;
output 	pc_out_25;
output 	pc_out_24;
output 	pc_out_27;
output 	pc_out_26;
input 	predicted_M;
input 	pc_plus_4_2;
input 	pc_plus_4_3;
input 	pc_plus_4_4;
input 	pc_plus_4_5;
input 	pc_plus_4_6;
input 	pc_plus_4_7;
input 	pc_plus_4_8;
input 	pc_plus_4_9;
input 	pc_plus_4_10;
input 	pc_plus_4_11;
input 	pc_plus_4_12;
input 	pc_plus_4_13;
input 	pc_plus_4_14;
input 	pc_plus_4_15;
input 	pc_plus_4_16;
input 	pc_plus_4_17;
input 	pc_plus_4_18;
input 	pc_plus_4_19;
input 	pc_plus_4_20;
input 	pc_plus_4_21;
input 	pc_plus_4_22;
input 	pc_plus_4_23;
input 	pc_plus_4_24;
input 	pc_plus_4_25;
input 	pc_plus_4_26;
input 	pc_plus_4_27;
output 	pc_out_1;
output 	pc_out_0;
output 	pc_out_29;
output 	pc_out_28;
output 	pc_out_31;
output 	pc_out_30;
input 	j_M;
input 	jal_M;
input 	branch_or_jump;
input 	branch_taken;
input 	jr_M;
input 	branch_or_jump1;
input 	predicted;
input 	pc_next;
input 	pc_next_1;
input 	pc_next_0;
input 	pc_next_3;
input 	pc_next_31;
input 	comb;
input 	pc_next_2;
input 	pc_next_21;
input 	pc_next_5;
input 	pc_next_51;
input 	pc_next_4;
input 	pc_next_41;
input 	pc_next_7;
input 	pc_next_71;
input 	pc_next_6;
input 	pc_next_61;
input 	pc_next_9;
input 	pc_next_91;
input 	pc_next_8;
input 	pc_next_81;
input 	pc_next_11;
input 	pc_next_111;
input 	pc_next_10;
input 	pc_next_101;
input 	pc_next_13;
input 	pc_next_131;
input 	pc_next_12;
input 	pc_next_121;
input 	pc_next_15;
input 	pc_next_151;
input 	pc_next_14;
input 	pc_next_141;
input 	pc_next_17;
input 	pc_next_171;
input 	pc_next_16;
input 	pc_next_161;
input 	pc_next_19;
input 	pc_next_191;
input 	pc_next_18;
input 	pc_next_181;
input 	pc_next_211;
input 	pc_next_212;
input 	pc_next_20;
input 	pc_next_201;
input 	pc_next_23;
input 	pc_next_231;
input 	pc_next_22;
input 	pc_next_221;
input 	pc_next_25;
input 	pc_next_251;
input 	pc_next_24;
input 	pc_next_241;
input 	pc_next_27;
input 	pc_next_271;
input 	pc_next_26;
input 	pc_next_261;
output 	pc_out_291;
output 	pc_out_292;
input 	pc_next_29;
input 	pc_next_28;
input 	pc_next_311;
input 	pc_next_30;
input 	comb1;
output 	pc_out_101;
input 	nRST;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \pc_out[3]~0_combout ;
wire \pc_out[2]~1_combout ;
wire \pc_out[5]~3_combout ;
wire \pc_out[4]~2_combout ;
wire \pc_out[7]~5_combout ;
wire \pc_out[6]~4_combout ;
wire \pc_out[9]~7_combout ;
wire \pc_out[8]~6_combout ;
wire \pc_out[11]~9_combout ;
wire \pc_out[10]~8_combout ;
wire \pc_out[13]~11_combout ;
wire \pc_out[12]~10_combout ;
wire \pc_out[15]~13_combout ;
wire \pc_out[14]~12_combout ;
wire \pc_out[17]~15_combout ;
wire \pc_out[16]~14_combout ;
wire \pc_out[19]~17_combout ;
wire \pc_out[18]~16_combout ;
wire \pc_out[21]~19_combout ;
wire \pc_out[20]~18_combout ;
wire \pc_out[23]~21_combout ;
wire \pc_out[22]~20_combout ;
wire \pc_out[25]~23_combout ;
wire \pc_out[24]~22_combout ;
wire \pc_out[27]~25_combout ;
wire \pc_out[26]~24_combout ;
wire \pc_out[1]~28_combout ;


// Location: FF_X56_Y37_N1
dffeas \pc_out[3] (
	.clk(CLK),
	.d(\pc_out[3]~0_combout ),
	.asdata(pc_next_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_3),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[3] .is_wysiwyg = "true";
defparam \pc_out[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N15
dffeas \pc_out[2] (
	.clk(CLK),
	.d(\pc_out[2]~1_combout ),
	.asdata(pc_next_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_2),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[2] .is_wysiwyg = "true";
defparam \pc_out[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N5
dffeas \pc_out[5] (
	.clk(CLK),
	.d(\pc_out[5]~3_combout ),
	.asdata(pc_next_51),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_5),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[5] .is_wysiwyg = "true";
defparam \pc_out[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N9
dffeas \pc_out[4] (
	.clk(CLK),
	.d(\pc_out[4]~2_combout ),
	.asdata(pc_next_41),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_4),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[4] .is_wysiwyg = "true";
defparam \pc_out[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N17
dffeas \pc_out[7] (
	.clk(CLK),
	.d(\pc_out[7]~5_combout ),
	.asdata(pc_next_71),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_7),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[7] .is_wysiwyg = "true";
defparam \pc_out[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N3
dffeas \pc_out[6] (
	.clk(CLK),
	.d(\pc_out[6]~4_combout ),
	.asdata(pc_next_61),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_6),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[6] .is_wysiwyg = "true";
defparam \pc_out[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N29
dffeas \pc_out[9] (
	.clk(CLK),
	.d(\pc_out[9]~7_combout ),
	.asdata(pc_next_91),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_9),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[9] .is_wysiwyg = "true";
defparam \pc_out[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N31
dffeas \pc_out[8] (
	.clk(CLK),
	.d(\pc_out[8]~6_combout ),
	.asdata(pc_next_81),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_8),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[8] .is_wysiwyg = "true";
defparam \pc_out[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N13
dffeas \pc_out[11] (
	.clk(CLK),
	.d(\pc_out[11]~9_combout ),
	.asdata(pc_next_111),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_11),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[11] .is_wysiwyg = "true";
defparam \pc_out[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N1
dffeas \pc_out[10] (
	.clk(CLK),
	.d(\pc_out[10]~8_combout ),
	.asdata(pc_next_101),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_10),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[10] .is_wysiwyg = "true";
defparam \pc_out[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N31
dffeas \pc_out[13] (
	.clk(CLK),
	.d(\pc_out[13]~11_combout ),
	.asdata(pc_next_131),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_13),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[13] .is_wysiwyg = "true";
defparam \pc_out[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N7
dffeas \pc_out[12] (
	.clk(CLK),
	.d(\pc_out[12]~10_combout ),
	.asdata(pc_next_121),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_12),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[12] .is_wysiwyg = "true";
defparam \pc_out[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N13
dffeas \pc_out[15] (
	.clk(CLK),
	.d(\pc_out[15]~13_combout ),
	.asdata(pc_next_151),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_15),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[15] .is_wysiwyg = "true";
defparam \pc_out[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N19
dffeas \pc_out[14] (
	.clk(CLK),
	.d(\pc_out[14]~12_combout ),
	.asdata(pc_next_141),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_14),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[14] .is_wysiwyg = "true";
defparam \pc_out[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N25
dffeas \pc_out[17] (
	.clk(CLK),
	.d(\pc_out[17]~15_combout ),
	.asdata(pc_next_171),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_17),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[17] .is_wysiwyg = "true";
defparam \pc_out[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y37_N5
dffeas \pc_out[16] (
	.clk(CLK),
	.d(\pc_out[16]~14_combout ),
	.asdata(pc_next_161),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_16),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[16] .is_wysiwyg = "true";
defparam \pc_out[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N9
dffeas \pc_out[19] (
	.clk(CLK),
	.d(\pc_out[19]~17_combout ),
	.asdata(pc_next_191),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_19),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[19] .is_wysiwyg = "true";
defparam \pc_out[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N23
dffeas \pc_out[18] (
	.clk(CLK),
	.d(\pc_out[18]~16_combout ),
	.asdata(pc_next_181),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_18),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[18] .is_wysiwyg = "true";
defparam \pc_out[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N11
dffeas \pc_out[21] (
	.clk(CLK),
	.d(\pc_out[21]~19_combout ),
	.asdata(pc_next_212),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_21),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[21] .is_wysiwyg = "true";
defparam \pc_out[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N7
dffeas \pc_out[20] (
	.clk(CLK),
	.d(\pc_out[20]~18_combout ),
	.asdata(pc_next_201),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_20),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[20] .is_wysiwyg = "true";
defparam \pc_out[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N13
dffeas \pc_out[23] (
	.clk(CLK),
	.d(\pc_out[23]~21_combout ),
	.asdata(pc_next_231),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_23),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[23] .is_wysiwyg = "true";
defparam \pc_out[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N7
dffeas \pc_out[22] (
	.clk(CLK),
	.d(\pc_out[22]~20_combout ),
	.asdata(pc_next_221),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_22),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[22] .is_wysiwyg = "true";
defparam \pc_out[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N29
dffeas \pc_out[25] (
	.clk(CLK),
	.d(\pc_out[25]~23_combout ),
	.asdata(pc_next_251),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_25),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[25] .is_wysiwyg = "true";
defparam \pc_out[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N31
dffeas \pc_out[24] (
	.clk(CLK),
	.d(\pc_out[24]~22_combout ),
	.asdata(pc_next_241),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_24),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[24] .is_wysiwyg = "true";
defparam \pc_out[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y39_N17
dffeas \pc_out[27] (
	.clk(CLK),
	.d(\pc_out[27]~25_combout ),
	.asdata(pc_next_271),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_27),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[27] .is_wysiwyg = "true";
defparam \pc_out[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N25
dffeas \pc_out[26] (
	.clk(CLK),
	.d(\pc_out[26]~24_combout ),
	.asdata(pc_next_261),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(pc_next),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_26),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[26] .is_wysiwyg = "true";
defparam \pc_out[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N29
dffeas \pc_out[1] (
	.clk(CLK),
	.d(pc_next_1),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_out[1]~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_1),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[1] .is_wysiwyg = "true";
defparam \pc_out[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N23
dffeas \pc_out[0] (
	.clk(CLK),
	.d(pc_next_0),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc_out[1]~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_0),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[0] .is_wysiwyg = "true";
defparam \pc_out[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N5
dffeas \pc_out[29] (
	.clk(CLK),
	.d(pc_next_29),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_29),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[29] .is_wysiwyg = "true";
defparam \pc_out[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N23
dffeas \pc_out[28] (
	.clk(CLK),
	.d(pc_next_28),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_28),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[28] .is_wysiwyg = "true";
defparam \pc_out[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N1
dffeas \pc_out[31] (
	.clk(CLK),
	.d(pc_next_311),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_31),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[31] .is_wysiwyg = "true";
defparam \pc_out[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N15
dffeas \pc_out[30] (
	.clk(CLK),
	.d(pc_next_30),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_out_30),
	.prn(vcc));
// synopsys translate_off
defparam \pc_out[30] .is_wysiwyg = "true";
defparam \pc_out[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N30
cycloneive_lcell_comb \pc_out[29]~29 (
// Equation(s):
// pc_out_291 = (\branch_or_jump~0_combout  & ((\jr_M~q ) # (\predicted_M~q  $ (!\branch_taken~0_combout ))))

	.dataa(jr_M),
	.datab(branch_or_jump),
	.datac(predicted_M),
	.datad(branch_taken),
	.cin(gnd),
	.combout(pc_out_291),
	.cout());
// synopsys translate_off
defparam \pc_out[29]~29 .lut_mask = 16'hC88C;
defparam \pc_out[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N16
cycloneive_lcell_comb \pc_out[29]~30 (
// Equation(s):
// pc_out_292 = (\branch_or_jump~0_combout  & ((\jr_M~q ) # ((!\predicted_M~q  & \branch_taken~0_combout ))))

	.dataa(jr_M),
	.datab(branch_or_jump),
	.datac(predicted_M),
	.datad(branch_taken),
	.cin(gnd),
	.combout(pc_out_292),
	.cout());
// synopsys translate_off
defparam \pc_out[29]~30 .lut_mask = 16'h8C88;
defparam \pc_out[29]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N6
cycloneive_lcell_comb \pc_out[10]~31 (
// Equation(s):
// pc_out_101 = (\jal_M~q ) # ((\j_M~q ) # ((!\jr_M~q  & \branch_taken~0_combout )))

	.dataa(jr_M),
	.datab(jal_M),
	.datac(j_M),
	.datad(branch_taken),
	.cin(gnd),
	.combout(pc_out_101),
	.cout());
// synopsys translate_off
defparam \pc_out[10]~31 .lut_mask = 16'hFDFC;
defparam \pc_out[10]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N0
cycloneive_lcell_comb \pc_out[3]~0 (
// Equation(s):
// \pc_out[3]~0_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[3]~2_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[3]~10_combout )))

	.dataa(pc_plus_4_3),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_3),
	.cin(gnd),
	.combout(\pc_out[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[3]~0 .lut_mask = 16'hBB88;
defparam \pc_out[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N14
cycloneive_lcell_comb \pc_out[2]~1 (
// Equation(s):
// \pc_out[2]~1_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[2]~0_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[2]~14_combout )))

	.dataa(pc_plus_4_2),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_2),
	.cin(gnd),
	.combout(\pc_out[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[2]~1 .lut_mask = 16'hBB88;
defparam \pc_out[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N4
cycloneive_lcell_comb \pc_out[5]~3 (
// Equation(s):
// \pc_out[5]~3_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[5]~6_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[5]~18_combout )))

	.dataa(branch_or_jump1),
	.datab(pc_plus_4_5),
	.datac(gnd),
	.datad(pc_next_5),
	.cin(gnd),
	.combout(\pc_out[5]~3_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[5]~3 .lut_mask = 16'hDD88;
defparam \pc_out[5]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N8
cycloneive_lcell_comb \pc_out[4]~2 (
// Equation(s):
// \pc_out[4]~2_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[4]~4_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[4]~22_combout )))

	.dataa(pc_plus_4_4),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_4),
	.cin(gnd),
	.combout(\pc_out[4]~2_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[4]~2 .lut_mask = 16'hBB88;
defparam \pc_out[4]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N16
cycloneive_lcell_comb \pc_out[7]~5 (
// Equation(s):
// \pc_out[7]~5_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[7]~10_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[7]~26_combout )))

	.dataa(branch_or_jump1),
	.datab(pc_plus_4_7),
	.datac(gnd),
	.datad(pc_next_7),
	.cin(gnd),
	.combout(\pc_out[7]~5_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[7]~5 .lut_mask = 16'hDD88;
defparam \pc_out[7]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N2
cycloneive_lcell_comb \pc_out[6]~4 (
// Equation(s):
// \pc_out[6]~4_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[6]~8_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[6]~30_combout )))

	.dataa(branch_or_jump1),
	.datab(pc_plus_4_6),
	.datac(gnd),
	.datad(pc_next_6),
	.cin(gnd),
	.combout(\pc_out[6]~4_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[6]~4 .lut_mask = 16'hDD88;
defparam \pc_out[6]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N28
cycloneive_lcell_comb \pc_out[9]~7 (
// Equation(s):
// \pc_out[9]~7_combout  = (\branch_or_jump~1_combout  & ((\pc_plus_4[9]~14_combout ))) # (!\branch_or_jump~1_combout  & (\pc_next[9]~34_combout ))

	.dataa(pc_next_9),
	.datab(pc_plus_4_9),
	.datac(gnd),
	.datad(branch_or_jump1),
	.cin(gnd),
	.combout(\pc_out[9]~7_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[9]~7 .lut_mask = 16'hCCAA;
defparam \pc_out[9]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N30
cycloneive_lcell_comb \pc_out[8]~6 (
// Equation(s):
// \pc_out[8]~6_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[8]~12_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[8]~38_combout )))

	.dataa(branch_or_jump1),
	.datab(pc_plus_4_8),
	.datac(gnd),
	.datad(pc_next_8),
	.cin(gnd),
	.combout(\pc_out[8]~6_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[8]~6 .lut_mask = 16'hDD88;
defparam \pc_out[8]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N12
cycloneive_lcell_comb \pc_out[11]~9 (
// Equation(s):
// \pc_out[11]~9_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[11]~18_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[11]~42_combout )))

	.dataa(branch_or_jump1),
	.datab(pc_plus_4_11),
	.datac(gnd),
	.datad(pc_next_11),
	.cin(gnd),
	.combout(\pc_out[11]~9_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[11]~9 .lut_mask = 16'hDD88;
defparam \pc_out[11]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N0
cycloneive_lcell_comb \pc_out[10]~8 (
// Equation(s):
// \pc_out[10]~8_combout  = (\branch_or_jump~1_combout  & ((\pc_plus_4[10]~16_combout ))) # (!\branch_or_jump~1_combout  & (\pc_next[10]~46_combout ))

	.dataa(pc_next_10),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_plus_4_10),
	.cin(gnd),
	.combout(\pc_out[10]~8_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[10]~8 .lut_mask = 16'hEE22;
defparam \pc_out[10]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N30
cycloneive_lcell_comb \pc_out[13]~11 (
// Equation(s):
// \pc_out[13]~11_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[13]~22_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[13]~50_combout )))

	.dataa(pc_plus_4_13),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_13),
	.cin(gnd),
	.combout(\pc_out[13]~11_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[13]~11 .lut_mask = 16'hBB88;
defparam \pc_out[13]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N6
cycloneive_lcell_comb \pc_out[12]~10 (
// Equation(s):
// \pc_out[12]~10_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[12]~20_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[12]~54_combout )))

	.dataa(pc_plus_4_12),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_12),
	.cin(gnd),
	.combout(\pc_out[12]~10_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[12]~10 .lut_mask = 16'hBB88;
defparam \pc_out[12]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N12
cycloneive_lcell_comb \pc_out[15]~13 (
// Equation(s):
// \pc_out[15]~13_combout  = (\branch_or_jump~1_combout  & ((\pc_plus_4[15]~26_combout ))) # (!\branch_or_jump~1_combout  & (\pc_next[15]~58_combout ))

	.dataa(pc_next_15),
	.datab(pc_plus_4_15),
	.datac(gnd),
	.datad(branch_or_jump1),
	.cin(gnd),
	.combout(\pc_out[15]~13_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[15]~13 .lut_mask = 16'hCCAA;
defparam \pc_out[15]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N18
cycloneive_lcell_comb \pc_out[14]~12 (
// Equation(s):
// \pc_out[14]~12_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[14]~24_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[14]~62_combout )))

	.dataa(pc_plus_4_14),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_14),
	.cin(gnd),
	.combout(\pc_out[14]~12_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[14]~12 .lut_mask = 16'hBB88;
defparam \pc_out[14]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N24
cycloneive_lcell_comb \pc_out[17]~15 (
// Equation(s):
// \pc_out[17]~15_combout  = (\branch_or_jump~1_combout  & ((\pc_plus_4[17]~30_combout ))) # (!\branch_or_jump~1_combout  & (\pc_next[17]~66_combout ))

	.dataa(pc_next_17),
	.datab(pc_plus_4_17),
	.datac(gnd),
	.datad(branch_or_jump1),
	.cin(gnd),
	.combout(\pc_out[17]~15_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[17]~15 .lut_mask = 16'hCCAA;
defparam \pc_out[17]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N4
cycloneive_lcell_comb \pc_out[16]~14 (
// Equation(s):
// \pc_out[16]~14_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[16]~28_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[16]~70_combout )))

	.dataa(pc_plus_4_16),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_16),
	.cin(gnd),
	.combout(\pc_out[16]~14_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[16]~14 .lut_mask = 16'hBB88;
defparam \pc_out[16]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N8
cycloneive_lcell_comb \pc_out[19]~17 (
// Equation(s):
// \pc_out[19]~17_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[19]~34_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[19]~74_combout )))

	.dataa(pc_plus_4_19),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_19),
	.cin(gnd),
	.combout(\pc_out[19]~17_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[19]~17 .lut_mask = 16'hBB88;
defparam \pc_out[19]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N22
cycloneive_lcell_comb \pc_out[18]~16 (
// Equation(s):
// \pc_out[18]~16_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[18]~32_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[18]~78_combout )))

	.dataa(pc_plus_4_18),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_18),
	.cin(gnd),
	.combout(\pc_out[18]~16_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[18]~16 .lut_mask = 16'hBB88;
defparam \pc_out[18]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N10
cycloneive_lcell_comb \pc_out[21]~19 (
// Equation(s):
// \pc_out[21]~19_combout  = (\branch_or_jump~1_combout  & ((\pc_plus_4[21]~38_combout ))) # (!\branch_or_jump~1_combout  & (\pc_next[21]~82_combout ))

	.dataa(pc_next_211),
	.datab(pc_plus_4_21),
	.datac(gnd),
	.datad(branch_or_jump1),
	.cin(gnd),
	.combout(\pc_out[21]~19_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[21]~19 .lut_mask = 16'hCCAA;
defparam \pc_out[21]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N6
cycloneive_lcell_comb \pc_out[20]~18 (
// Equation(s):
// \pc_out[20]~18_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[20]~36_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[20]~86_combout )))

	.dataa(pc_plus_4_20),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_20),
	.cin(gnd),
	.combout(\pc_out[20]~18_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[20]~18 .lut_mask = 16'hBB88;
defparam \pc_out[20]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N12
cycloneive_lcell_comb \pc_out[23]~21 (
// Equation(s):
// \pc_out[23]~21_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[23]~42_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[23]~90_combout )))

	.dataa(branch_or_jump1),
	.datab(pc_plus_4_23),
	.datac(gnd),
	.datad(pc_next_23),
	.cin(gnd),
	.combout(\pc_out[23]~21_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[23]~21 .lut_mask = 16'hDD88;
defparam \pc_out[23]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N6
cycloneive_lcell_comb \pc_out[22]~20 (
// Equation(s):
// \pc_out[22]~20_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[22]~40_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[22]~94_combout )))

	.dataa(pc_plus_4_22),
	.datab(pc_next_22),
	.datac(gnd),
	.datad(branch_or_jump1),
	.cin(gnd),
	.combout(\pc_out[22]~20_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[22]~20 .lut_mask = 16'hAACC;
defparam \pc_out[22]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N28
cycloneive_lcell_comb \pc_out[25]~23 (
// Equation(s):
// \pc_out[25]~23_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[25]~46_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[25]~98_combout )))

	.dataa(branch_or_jump1),
	.datab(pc_plus_4_25),
	.datac(gnd),
	.datad(pc_next_25),
	.cin(gnd),
	.combout(\pc_out[25]~23_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[25]~23 .lut_mask = 16'hDD88;
defparam \pc_out[25]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N30
cycloneive_lcell_comb \pc_out[24]~22 (
// Equation(s):
// \pc_out[24]~22_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[24]~44_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[24]~102_combout )))

	.dataa(pc_plus_4_24),
	.datab(pc_next_24),
	.datac(gnd),
	.datad(branch_or_jump1),
	.cin(gnd),
	.combout(\pc_out[24]~22_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[24]~22 .lut_mask = 16'hAACC;
defparam \pc_out[24]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N16
cycloneive_lcell_comb \pc_out[27]~25 (
// Equation(s):
// \pc_out[27]~25_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[27]~50_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[27]~106_combout )))

	.dataa(pc_plus_4_27),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_27),
	.cin(gnd),
	.combout(\pc_out[27]~25_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[27]~25 .lut_mask = 16'hBB88;
defparam \pc_out[27]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N24
cycloneive_lcell_comb \pc_out[26]~24 (
// Equation(s):
// \pc_out[26]~24_combout  = (\branch_or_jump~1_combout  & (\pc_plus_4[26]~48_combout )) # (!\branch_or_jump~1_combout  & ((\pc_next[26]~110_combout )))

	.dataa(pc_plus_4_26),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(pc_next_26),
	.cin(gnd),
	.combout(\pc_out[26]~24_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[26]~24 .lut_mask = 16'hBB88;
defparam \pc_out[26]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N24
cycloneive_lcell_comb \pc_out[1]~28 (
// Equation(s):
// \pc_out[1]~28_combout  = ((predicted & \comb~3_combout )) # (!\branch_or_jump~1_combout )

	.dataa(predicted),
	.datab(branch_or_jump1),
	.datac(gnd),
	.datad(comb1),
	.cin(gnd),
	.combout(\pc_out[1]~28_combout ),
	.cout());
// synopsys translate_off
defparam \pc_out[1]~28 .lut_mask = 16'hBB33;
defparam \pc_out[1]~28 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module register_file (
	wsel_WB_1,
	wsel_WB_0,
	wsel_WB_3,
	wsel_WB_2,
	wsel_WB_4,
	regWrite_WB,
	wdat_WB_31,
	wdat_WB_30,
	wdat_WB_29,
	wdat_WB_28,
	wdat_WB_27,
	wdat_WB_26,
	wdat_WB_25,
	wdat_WB_24,
	wdat_WB_23,
	wdat_WB_22,
	wdat_WB_21,
	wdat_WB_20,
	wdat_WB_19,
	wdat_WB_18,
	wdat_WB_17,
	wdat_WB_16,
	wdat_WB_15,
	wdat_WB_14,
	wdat_WB_13,
	wdat_WB_12,
	wdat_WB_9,
	wdat_WB_8,
	wdat_WB_11,
	wdat_WB_10,
	wdat_WB_7,
	wdat_WB_6,
	wdat_WB_5,
	wdat_WB_2,
	wdat_WB_1,
	wdat_WB_0,
	wdat_WB_4,
	wdat_WB_3,
	instruction_D_16,
	instruction_D_17,
	instruction_D_18,
	instruction_D_19,
	instruction_D_22,
	instruction_D_21,
	instruction_D_24,
	instruction_D_23,
	Mux32,
	Mux321,
	Mux33,
	Mux331,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux36,
	Mux361,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux41,
	Mux411,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux44,
	Mux441,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux48,
	Mux481,
	Mux49,
	Mux491,
	Mux50,
	Mux501,
	Mux51,
	Mux511,
	Mux54,
	Mux541,
	Mux55,
	Mux551,
	Mux52,
	Mux521,
	Mux53,
	Mux531,
	Mux56,
	Mux561,
	Mux57,
	Mux571,
	Mux58,
	Mux581,
	Mux29,
	Mux291,
	Mux30,
	Mux301,
	Mux63,
	Mux631,
	Mux62,
	Mux621,
	Mux27,
	Mux271,
	Mux28,
	Mux281,
	Mux61,
	Mux611,
	Mux23,
	Mux231,
	Mux24,
	Mux241,
	Mux25,
	Mux251,
	Mux26,
	Mux261,
	Mux60,
	Mux601,
	Mux15,
	Mux151,
	Mux16,
	Mux161,
	Mux17,
	Mux171,
	Mux18,
	Mux181,
	Mux19,
	Mux191,
	Mux20,
	Mux201,
	Mux21,
	Mux211,
	Mux22,
	Mux221,
	Mux59,
	Mux591,
	Mux0,
	Mux01,
	Mux2,
	Mux210,
	Mux1,
	Mux11,
	Mux3,
	Mux31,
	Mux4,
	Mux410,
	Mux5,
	Mux510,
	Mux6,
	Mux64,
	Mux7,
	Mux71,
	Mux8,
	Mux81,
	Mux9,
	Mux91,
	Mux10,
	Mux101,
	Mux111,
	Mux112,
	Mux12,
	Mux121,
	Mux13,
	Mux131,
	Mux14,
	Mux141,
	Mux311,
	Mux312,
	nRST,
	CLK,
	devpor,
	devclrn,
	devoe);
input 	wsel_WB_1;
input 	wsel_WB_0;
input 	wsel_WB_3;
input 	wsel_WB_2;
input 	wsel_WB_4;
input 	regWrite_WB;
input 	wdat_WB_31;
input 	wdat_WB_30;
input 	wdat_WB_29;
input 	wdat_WB_28;
input 	wdat_WB_27;
input 	wdat_WB_26;
input 	wdat_WB_25;
input 	wdat_WB_24;
input 	wdat_WB_23;
input 	wdat_WB_22;
input 	wdat_WB_21;
input 	wdat_WB_20;
input 	wdat_WB_19;
input 	wdat_WB_18;
input 	wdat_WB_17;
input 	wdat_WB_16;
input 	wdat_WB_15;
input 	wdat_WB_14;
input 	wdat_WB_13;
input 	wdat_WB_12;
input 	wdat_WB_9;
input 	wdat_WB_8;
input 	wdat_WB_11;
input 	wdat_WB_10;
input 	wdat_WB_7;
input 	wdat_WB_6;
input 	wdat_WB_5;
input 	wdat_WB_2;
input 	wdat_WB_1;
input 	wdat_WB_0;
input 	wdat_WB_4;
input 	wdat_WB_3;
input 	instruction_D_16;
input 	instruction_D_17;
input 	instruction_D_18;
input 	instruction_D_19;
input 	instruction_D_22;
input 	instruction_D_21;
input 	instruction_D_24;
input 	instruction_D_23;
output 	Mux32;
output 	Mux321;
output 	Mux33;
output 	Mux331;
output 	Mux34;
output 	Mux341;
output 	Mux35;
output 	Mux351;
output 	Mux36;
output 	Mux361;
output 	Mux37;
output 	Mux371;
output 	Mux38;
output 	Mux381;
output 	Mux39;
output 	Mux391;
output 	Mux40;
output 	Mux401;
output 	Mux41;
output 	Mux411;
output 	Mux42;
output 	Mux421;
output 	Mux43;
output 	Mux431;
output 	Mux44;
output 	Mux441;
output 	Mux45;
output 	Mux451;
output 	Mux46;
output 	Mux461;
output 	Mux47;
output 	Mux471;
output 	Mux48;
output 	Mux481;
output 	Mux49;
output 	Mux491;
output 	Mux50;
output 	Mux501;
output 	Mux51;
output 	Mux511;
output 	Mux54;
output 	Mux541;
output 	Mux55;
output 	Mux551;
output 	Mux52;
output 	Mux521;
output 	Mux53;
output 	Mux531;
output 	Mux56;
output 	Mux561;
output 	Mux57;
output 	Mux571;
output 	Mux58;
output 	Mux581;
output 	Mux29;
output 	Mux291;
output 	Mux30;
output 	Mux301;
output 	Mux63;
output 	Mux631;
output 	Mux62;
output 	Mux621;
output 	Mux27;
output 	Mux271;
output 	Mux28;
output 	Mux281;
output 	Mux61;
output 	Mux611;
output 	Mux23;
output 	Mux231;
output 	Mux24;
output 	Mux241;
output 	Mux25;
output 	Mux251;
output 	Mux26;
output 	Mux261;
output 	Mux60;
output 	Mux601;
output 	Mux15;
output 	Mux151;
output 	Mux16;
output 	Mux161;
output 	Mux17;
output 	Mux171;
output 	Mux18;
output 	Mux181;
output 	Mux19;
output 	Mux191;
output 	Mux20;
output 	Mux201;
output 	Mux21;
output 	Mux211;
output 	Mux22;
output 	Mux221;
output 	Mux59;
output 	Mux591;
output 	Mux0;
output 	Mux01;
output 	Mux2;
output 	Mux210;
output 	Mux1;
output 	Mux11;
output 	Mux3;
output 	Mux31;
output 	Mux4;
output 	Mux410;
output 	Mux5;
output 	Mux510;
output 	Mux6;
output 	Mux64;
output 	Mux7;
output 	Mux71;
output 	Mux8;
output 	Mux81;
output 	Mux9;
output 	Mux91;
output 	Mux10;
output 	Mux101;
output 	Mux111;
output 	Mux112;
output 	Mux12;
output 	Mux121;
output 	Mux13;
output 	Mux131;
output 	Mux14;
output 	Mux141;
output 	Mux311;
output 	Mux312;
input 	nRST;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Mux32~2_combout ;
wire \Mux33~2_combout ;
wire \rfile[28][30]~q ;
wire \Mux34~4_combout ;
wire \rfile[7][27]~q ;
wire \Mux37~4_combout ;
wire \Mux38~2_combout ;
wire \rfile[16][24]~q ;
wire \Mux39~4_combout ;
wire \rfile[9][24]~q ;
wire \rfile[28][22]~q ;
wire \Mux44~12_combout ;
wire \rfile[5][18]~q ;
wire \Mux47~2_combout ;
wire \rfile[24][16]~q ;
wire \Mux51~12_combout ;
wire \Mux54~12_combout ;
wire \rfile[2][9]~q ;
wire \rfile[28][8]~q ;
wire \rfile[6][7]~q ;
wire \rfile[26][1]~q ;
wire \rfile[18][1]~q ;
wire \Mux30~2_combout ;
wire \rfile[4][1]~q ;
wire \Mux30~12_combout ;
wire \rfile[2][1]~q ;
wire \rfile[12][1]~q ;
wire \Mux62~2_combout ;
wire \Mux24~4_combout ;
wire \Mux25~2_combout ;
wire \Mux21~4_combout ;
wire \Mux21~12_combout ;
wire \Mux0~14_combout ;
wire \Mux7~2_combout ;
wire \Mux14~2_combout ;
wire \rfile[28][30]~feeder_combout ;
wire \rfile[7][27]~feeder_combout ;
wire \rfile[9][24]~feeder_combout ;
wire \rfile[28][22]~feeder_combout ;
wire \rfile[5][18]~feeder_combout ;
wire \rfile[24][16]~feeder_combout ;
wire \rfile[2][9]~feeder_combout ;
wire \rfile[28][8]~feeder_combout ;
wire \rfile[6][7]~feeder_combout ;
wire \rfile[2][1]~feeder_combout ;
wire \rfile[12][1]~feeder_combout ;
wire \Decoder0~2_combout ;
wire \Decoder0~4_combout ;
wire \rfile[17][31]~q ;
wire \Decoder0~3_combout ;
wire \rfile[21][31]~q ;
wire \Mux32~0_combout ;
wire \rfile[25][31]~feeder_combout ;
wire \Decoder0~0_combout ;
wire \Decoder0~1_combout ;
wire \rfile[25][31]~q ;
wire \Decoder0~5_combout ;
wire \rfile[29][31]~q ;
wire \Mux32~1_combout ;
wire \Decoder0~8_combout ;
wire \Decoder0~16_combout ;
wire \rfile[27][31]~q ;
wire \Decoder0~6_combout ;
wire \Decoder0~17_combout ;
wire \rfile[23][31]~q ;
wire \rfile[19][31]~feeder_combout ;
wire \Decoder0~18_combout ;
wire \rfile[19][31]~q ;
wire \Mux32~7_combout ;
wire \rfile[31][31]~feeder_combout ;
wire \Decoder0~19_combout ;
wire \rfile[31][31]~q ;
wire \Mux32~8_combout ;
wire \rfile[28][31]~feeder_combout ;
wire \Decoder0~15_combout ;
wire \rfile[28][31]~q ;
wire \Decoder0~13_combout ;
wire \rfile[24][31]~q ;
wire \Decoder0~14_combout ;
wire \rfile[16][31]~q ;
wire \Mux32~4_combout ;
wire \Mux32~5_combout ;
wire \Decoder0~7_combout ;
wire \rfile[22][31]~q ;
wire \Decoder0~11_combout ;
wire \rfile[30][31]~q ;
wire \Mux32~3_combout ;
wire \Mux32~6_combout ;
wire \rfile[11][31]~feeder_combout ;
wire \Decoder0~22_combout ;
wire \Decoder0~25_combout ;
wire \rfile[11][31]~q ;
wire \Decoder0~23_combout ;
wire \rfile[10][31]~q ;
wire \Mux32~10_combout ;
wire \rfile[9][31]~feeder_combout ;
wire \Decoder0~20_combout ;
wire \Decoder0~21_combout ;
wire \rfile[9][31]~q ;
wire \Mux32~11_combout ;
wire \Decoder0~26_combout ;
wire \Decoder0~27_combout ;
wire \rfile[6][31]~q ;
wire \Decoder0~28_combout ;
wire \Decoder0~29_combout ;
wire \rfile[5][31]~q ;
wire \Mux32~12_combout ;
wire \Mux32~13_combout ;
wire \Decoder0~34_combout ;
wire \rfile[2][31]~q ;
wire \Decoder0~32_combout ;
wire \rfile[3][31]~q ;
wire \Decoder0~33_combout ;
wire \rfile[1][31]~q ;
wire \Mux32~14_combout ;
wire \Mux32~15_combout ;
wire \Mux32~16_combout ;
wire \rfile[14][31]~feeder_combout ;
wire \Decoder0~35_combout ;
wire \rfile[14][31]~q ;
wire \Decoder0~38_combout ;
wire \rfile[15][31]~q ;
wire \Decoder0~37_combout ;
wire \rfile[12][31]~q ;
wire \Decoder0~36_combout ;
wire \rfile[13][31]~q ;
wire \Mux32~17_combout ;
wire \Mux32~18_combout ;
wire \rfile[21][30]~q ;
wire \rfile[29][30]~q ;
wire \rfile[25][30]~q ;
wire \rfile[17][30]~q ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \rfile[31][30]~q ;
wire \rfile[23][30]~q ;
wire \rfile[19][30]~q ;
wire \rfile[27][30]~q ;
wire \Mux33~7_combout ;
wire \Mux33~8_combout ;
wire \Decoder0~9_combout ;
wire \rfile[26][30]~q ;
wire \rfile[30][30]~q ;
wire \Mux33~3_combout ;
wire \rfile[24][30]~q ;
wire \Decoder0~12_combout ;
wire \rfile[20][30]~q ;
wire \rfile[16][30]~q ;
wire \Mux33~4_combout ;
wire \Mux33~5_combout ;
wire \Mux33~6_combout ;
wire \rfile[14][30]~q ;
wire \rfile[15][30]~q ;
wire \rfile[13][30]~q ;
wire \rfile[12][30]~q ;
wire \Mux33~17_combout ;
wire \Mux33~18_combout ;
wire \rfile[2][30]~feeder_combout ;
wire \rfile[2][30]~q ;
wire \rfile[3][30]~q ;
wire \rfile[1][30]~q ;
wire \Mux33~14_combout ;
wire \Mux33~15_combout ;
wire \rfile[9][30]~q ;
wire \Decoder0~24_combout ;
wire \rfile[8][30]~q ;
wire \rfile[10][30]~q ;
wire \Mux33~12_combout ;
wire \Mux33~13_combout ;
wire \Mux33~16_combout ;
wire \rfile[5][30]~q ;
wire \Mux33~10_combout ;
wire \rfile[6][30]~q ;
wire \Decoder0~31_combout ;
wire \rfile[7][30]~q ;
wire \Mux33~11_combout ;
wire \rfile[29][29]~q ;
wire \rfile[25][29]~feeder_combout ;
wire \rfile[25][29]~q ;
wire \rfile[21][29]~q ;
wire \rfile[17][29]~q ;
wire \Mux34~0_combout ;
wire \Mux34~1_combout ;
wire \rfile[20][29]~q ;
wire \rfile[28][29]~feeder_combout ;
wire \rfile[28][29]~q ;
wire \Mux34~5_combout ;
wire \rfile[30][29]~q ;
wire \rfile[22][29]~q ;
wire \rfile[18][29]~feeder_combout ;
wire \Decoder0~10_combout ;
wire \rfile[18][29]~q ;
wire \rfile[26][29]~feeder_combout ;
wire \rfile[26][29]~q ;
wire \Mux34~2_combout ;
wire \Mux34~3_combout ;
wire \Mux34~6_combout ;
wire \rfile[31][29]~q ;
wire \rfile[23][29]~q ;
wire \rfile[19][29]~q ;
wire \Mux34~7_combout ;
wire \rfile[27][29]~q ;
wire \Mux34~8_combout ;
wire \rfile[11][29]~q ;
wire \rfile[9][29]~q ;
wire \rfile[10][29]~q ;
wire \rfile[8][29]~q ;
wire \Mux34~10_combout ;
wire \Mux34~11_combout ;
wire \rfile[13][29]~q ;
wire \rfile[12][29]~q ;
wire \Mux34~17_combout ;
wire \rfile[15][29]~q ;
wire \rfile[14][29]~q ;
wire \Mux34~18_combout ;
wire \rfile[6][29]~q ;
wire \Decoder0~30_combout ;
wire \rfile[4][29]~q ;
wire \rfile[5][29]~q ;
wire \Mux34~12_combout ;
wire \Mux34~13_combout ;
wire \rfile[2][29]~q ;
wire \rfile[3][29]~q ;
wire \rfile[1][29]~feeder_combout ;
wire \rfile[1][29]~q ;
wire \Mux34~14_combout ;
wire \Mux34~15_combout ;
wire \Mux34~16_combout ;
wire \rfile[31][28]~q ;
wire \rfile[23][28]~q ;
wire \rfile[27][28]~q ;
wire \rfile[19][28]~q ;
wire \Mux35~7_combout ;
wire \Mux35~8_combout ;
wire \rfile[24][28]~q ;
wire \rfile[16][28]~q ;
wire \rfile[20][28]~q ;
wire \Mux35~4_combout ;
wire \Mux35~5_combout ;
wire \rfile[26][28]~q ;
wire \rfile[30][28]~q ;
wire \rfile[18][28]~q ;
wire \rfile[22][28]~q ;
wire \Mux35~2_combout ;
wire \Mux35~3_combout ;
wire \Mux35~6_combout ;
wire \rfile[21][28]~q ;
wire \rfile[29][28]~q ;
wire \rfile[17][28]~q ;
wire \rfile[25][28]~q ;
wire \Mux35~0_combout ;
wire \Mux35~1_combout ;
wire \rfile[14][28]~feeder_combout ;
wire \rfile[14][28]~q ;
wire \rfile[15][28]~q ;
wire \rfile[13][28]~q ;
wire \rfile[12][28]~q ;
wire \Mux35~17_combout ;
wire \Mux35~18_combout ;
wire \rfile[3][28]~q ;
wire \rfile[1][28]~q ;
wire \Mux35~14_combout ;
wire \rfile[2][28]~q ;
wire \Mux35~15_combout ;
wire \rfile[11][28]~feeder_combout ;
wire \rfile[11][28]~q ;
wire \rfile[9][28]~q ;
wire \rfile[8][28]~q ;
wire \rfile[10][28]~q ;
wire \Mux35~12_combout ;
wire \Mux35~13_combout ;
wire \Mux35~16_combout ;
wire \rfile[4][28]~q ;
wire \rfile[5][28]~q ;
wire \Mux35~10_combout ;
wire \rfile[7][28]~q ;
wire \rfile[6][28]~q ;
wire \Mux35~11_combout ;
wire \rfile[31][27]~q ;
wire \rfile[27][27]~q ;
wire \rfile[23][27]~q ;
wire \Mux36~7_combout ;
wire \Mux36~8_combout ;
wire \rfile[25][27]~feeder_combout ;
wire \rfile[25][27]~q ;
wire \rfile[29][27]~q ;
wire \rfile[17][27]~q ;
wire \rfile[21][27]~q ;
wire \Mux36~0_combout ;
wire \Mux36~1_combout ;
wire \rfile[30][27]~q ;
wire \rfile[26][27]~q ;
wire \rfile[18][27]~q ;
wire \Mux36~2_combout ;
wire \Mux36~3_combout ;
wire \rfile[24][27]~q ;
wire \rfile[16][27]~q ;
wire \Mux36~4_combout ;
wire \rfile[20][27]~feeder_combout ;
wire \rfile[20][27]~q ;
wire \Mux36~5_combout ;
wire \Mux36~6_combout ;
wire \rfile[13][27]~q ;
wire \rfile[12][27]~q ;
wire \Mux36~17_combout ;
wire \rfile[14][27]~q ;
wire \rfile[15][27]~q ;
wire \Mux36~18_combout ;
wire \rfile[6][27]~q ;
wire \rfile[5][27]~q ;
wire \rfile[4][27]~q ;
wire \Mux36~12_combout ;
wire \Mux36~13_combout ;
wire \rfile[2][27]~q ;
wire \rfile[1][27]~q ;
wire \rfile[3][27]~q ;
wire \Mux36~14_combout ;
wire \Mux36~15_combout ;
wire \Mux36~16_combout ;
wire \rfile[11][27]~feeder_combout ;
wire \rfile[11][27]~q ;
wire \rfile[8][27]~q ;
wire \rfile[10][27]~q ;
wire \Mux36~10_combout ;
wire \rfile[9][27]~q ;
wire \Mux36~11_combout ;
wire \rfile[31][26]~feeder_combout ;
wire \rfile[31][26]~q ;
wire \rfile[23][26]~q ;
wire \rfile[27][26]~q ;
wire \rfile[19][26]~q ;
wire \Mux37~7_combout ;
wire \Mux37~8_combout ;
wire \rfile[24][26]~q ;
wire \rfile[28][26]~q ;
wire \Mux37~5_combout ;
wire \rfile[22][26]~q ;
wire \Mux37~2_combout ;
wire \rfile[26][26]~q ;
wire \rfile[30][26]~q ;
wire \Mux37~3_combout ;
wire \Mux37~6_combout ;
wire \rfile[29][26]~feeder_combout ;
wire \rfile[29][26]~q ;
wire \rfile[21][26]~feeder_combout ;
wire \rfile[21][26]~q ;
wire \rfile[25][26]~q ;
wire \Mux37~0_combout ;
wire \Mux37~1_combout ;
wire \rfile[9][26]~feeder_combout ;
wire \rfile[9][26]~q ;
wire \rfile[8][26]~q ;
wire \Mux37~12_combout ;
wire \Mux37~13_combout ;
wire \rfile[2][26]~feeder_combout ;
wire \rfile[2][26]~q ;
wire \rfile[3][26]~q ;
wire \rfile[1][26]~q ;
wire \Mux37~14_combout ;
wire \Mux37~15_combout ;
wire \Mux37~16_combout ;
wire \rfile[4][26]~q ;
wire \rfile[5][26]~q ;
wire \Mux37~10_combout ;
wire \rfile[7][26]~q ;
wire \rfile[6][26]~q ;
wire \Mux37~11_combout ;
wire \rfile[12][26]~q ;
wire \rfile[13][26]~q ;
wire \Mux37~17_combout ;
wire \rfile[14][26]~q ;
wire \rfile[15][26]~q ;
wire \Mux37~18_combout ;
wire \rfile[23][25]~q ;
wire \Mux38~7_combout ;
wire \rfile[31][25]~q ;
wire \rfile[27][25]~q ;
wire \Mux38~8_combout ;
wire \rfile[29][25]~q ;
wire \rfile[25][25]~q ;
wire \rfile[17][25]~q ;
wire \rfile[21][25]~feeder_combout ;
wire \rfile[21][25]~q ;
wire \Mux38~0_combout ;
wire \Mux38~1_combout ;
wire \rfile[22][25]~q ;
wire \rfile[30][25]~feeder_combout ;
wire \rfile[30][25]~q ;
wire \Mux38~3_combout ;
wire \rfile[20][25]~q ;
wire \rfile[16][25]~q ;
wire \rfile[24][25]~feeder_combout ;
wire \rfile[24][25]~q ;
wire \Mux38~4_combout ;
wire \Mux38~5_combout ;
wire \Mux38~6_combout ;
wire \rfile[14][25]~q ;
wire \rfile[15][25]~q ;
wire \rfile[12][25]~q ;
wire \rfile[13][25]~q ;
wire \Mux38~17_combout ;
wire \Mux38~18_combout ;
wire \rfile[11][25]~feeder_combout ;
wire \rfile[11][25]~q ;
wire \rfile[9][25]~q ;
wire \rfile[10][25]~q ;
wire \rfile[8][25]~q ;
wire \Mux38~10_combout ;
wire \Mux38~11_combout ;
wire \rfile[7][25]~q ;
wire \rfile[6][25]~q ;
wire \rfile[5][25]~q ;
wire \rfile[4][25]~q ;
wire \Mux38~12_combout ;
wire \Mux38~13_combout ;
wire \rfile[3][25]~q ;
wire \rfile[1][25]~q ;
wire \Mux38~14_combout ;
wire \rfile[2][25]~feeder_combout ;
wire \rfile[2][25]~q ;
wire \Mux38~15_combout ;
wire \Mux38~16_combout ;
wire \rfile[29][24]~q ;
wire \rfile[21][24]~q ;
wire \rfile[25][24]~q ;
wire \rfile[17][24]~q ;
wire \Mux39~0_combout ;
wire \Mux39~1_combout ;
wire \rfile[18][24]~q ;
wire \rfile[22][24]~q ;
wire \Mux39~2_combout ;
wire \rfile[30][24]~q ;
wire \rfile[26][24]~q ;
wire \Mux39~3_combout ;
wire \rfile[28][24]~q ;
wire \rfile[24][24]~q ;
wire \Mux39~5_combout ;
wire \Mux39~6_combout ;
wire \rfile[23][24]~feeder_combout ;
wire \rfile[23][24]~q ;
wire \rfile[31][24]~q ;
wire \rfile[27][24]~q ;
wire \rfile[19][24]~q ;
wire \Mux39~7_combout ;
wire \Mux39~8_combout ;
wire \rfile[7][24]~q ;
wire \rfile[6][24]~feeder_combout ;
wire \rfile[6][24]~q ;
wire \rfile[5][24]~q ;
wire \Mux39~10_combout ;
wire \Mux39~11_combout ;
wire \rfile[2][24]~feeder_combout ;
wire \rfile[2][24]~q ;
wire \rfile[1][24]~q ;
wire \rfile[3][24]~q ;
wire \Mux39~14_combout ;
wire \Mux39~15_combout ;
wire \rfile[11][24]~feeder_combout ;
wire \rfile[11][24]~q ;
wire \rfile[8][24]~q ;
wire \rfile[10][24]~q ;
wire \Mux39~12_combout ;
wire \Mux39~13_combout ;
wire \Mux39~16_combout ;
wire \rfile[15][24]~feeder_combout ;
wire \rfile[15][24]~q ;
wire \rfile[14][24]~q ;
wire \rfile[12][24]~q ;
wire \rfile[13][24]~feeder_combout ;
wire \rfile[13][24]~q ;
wire \Mux39~17_combout ;
wire \Mux39~18_combout ;
wire \rfile[25][23]~feeder_combout ;
wire \rfile[25][23]~q ;
wire \rfile[29][23]~q ;
wire \rfile[21][23]~q ;
wire \rfile[17][23]~feeder_combout ;
wire \rfile[17][23]~q ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \rfile[27][23]~q ;
wire \rfile[31][23]~q ;
wire \rfile[19][23]~q ;
wire \rfile[23][23]~q ;
wire \Mux40~7_combout ;
wire \Mux40~8_combout ;
wire \rfile[20][23]~feeder_combout ;
wire \rfile[20][23]~q ;
wire \rfile[28][23]~q ;
wire \rfile[16][23]~q ;
wire \rfile[24][23]~q ;
wire \Mux40~4_combout ;
wire \Mux40~5_combout ;
wire \rfile[22][23]~feeder_combout ;
wire \rfile[22][23]~q ;
wire \rfile[30][23]~q ;
wire \rfile[18][23]~q ;
wire \rfile[26][23]~feeder_combout ;
wire \rfile[26][23]~q ;
wire \Mux40~2_combout ;
wire \Mux40~3_combout ;
wire \Mux40~6_combout ;
wire \rfile[2][23]~feeder_combout ;
wire \rfile[2][23]~q ;
wire \rfile[3][23]~q ;
wire \rfile[1][23]~q ;
wire \Mux40~14_combout ;
wire \Mux40~15_combout ;
wire \rfile[7][23]~q ;
wire \rfile[5][23]~q ;
wire \rfile[4][23]~q ;
wire \Mux40~12_combout ;
wire \Mux40~13_combout ;
wire \Mux40~16_combout ;
wire \rfile[11][23]~q ;
wire \rfile[9][23]~q ;
wire \rfile[8][23]~q ;
wire \rfile[10][23]~q ;
wire \Mux40~10_combout ;
wire \Mux40~11_combout ;
wire \rfile[13][23]~q ;
wire \rfile[12][23]~q ;
wire \Mux40~17_combout ;
wire \rfile[14][23]~q ;
wire \rfile[15][23]~feeder_combout ;
wire \rfile[15][23]~q ;
wire \Mux40~18_combout ;
wire \rfile[29][22]~feeder_combout ;
wire \rfile[29][22]~q ;
wire \rfile[21][22]~q ;
wire \rfile[17][22]~q ;
wire \rfile[25][22]~q ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \rfile[19][22]~q ;
wire \rfile[27][22]~q ;
wire \Mux41~7_combout ;
wire \rfile[31][22]~q ;
wire \rfile[23][22]~q ;
wire \Mux41~8_combout ;
wire \rfile[24][22]~feeder_combout ;
wire \rfile[24][22]~q ;
wire \rfile[16][22]~q ;
wire \rfile[20][22]~q ;
wire \Mux41~4_combout ;
wire \Mux41~5_combout ;
wire \rfile[30][22]~q ;
wire \rfile[26][22]~q ;
wire \rfile[22][22]~q ;
wire \rfile[18][22]~q ;
wire \Mux41~2_combout ;
wire \Mux41~3_combout ;
wire \Mux41~6_combout ;
wire \rfile[14][22]~feeder_combout ;
wire \rfile[14][22]~q ;
wire \rfile[13][22]~q ;
wire \rfile[12][22]~q ;
wire \Mux41~17_combout ;
wire \rfile[15][22]~feeder_combout ;
wire \rfile[15][22]~q ;
wire \Mux41~18_combout ;
wire \rfile[2][22]~q ;
wire \rfile[1][22]~q ;
wire \rfile[3][22]~q ;
wire \Mux41~14_combout ;
wire \Mux41~15_combout ;
wire \rfile[11][22]~feeder_combout ;
wire \rfile[11][22]~q ;
wire \rfile[9][22]~q ;
wire \rfile[8][22]~q ;
wire \rfile[10][22]~q ;
wire \Mux41~12_combout ;
wire \Mux41~13_combout ;
wire \Mux41~16_combout ;
wire \rfile[6][22]~feeder_combout ;
wire \rfile[6][22]~q ;
wire \rfile[7][22]~q ;
wire \rfile[4][22]~q ;
wire \rfile[5][22]~q ;
wire \Mux41~10_combout ;
wire \Mux41~11_combout ;
wire \rfile[29][21]~q ;
wire \rfile[25][21]~q ;
wire \rfile[21][21]~q ;
wire \rfile[17][21]~q ;
wire \Mux42~0_combout ;
wire \Mux42~1_combout ;
wire \rfile[27][21]~q ;
wire \rfile[31][21]~q ;
wire \rfile[19][21]~q ;
wire \rfile[23][21]~q ;
wire \Mux42~7_combout ;
wire \Mux42~8_combout ;
wire \rfile[24][21]~q ;
wire \rfile[16][21]~q ;
wire \Mux42~4_combout ;
wire \rfile[28][21]~q ;
wire \Mux42~5_combout ;
wire \rfile[30][21]~q ;
wire \rfile[22][21]~q ;
wire \rfile[26][21]~feeder_combout ;
wire \rfile[26][21]~q ;
wire \rfile[18][21]~feeder_combout ;
wire \rfile[18][21]~q ;
wire \Mux42~2_combout ;
wire \Mux42~3_combout ;
wire \Mux42~6_combout ;
wire \rfile[14][21]~feeder_combout ;
wire \rfile[14][21]~q ;
wire \rfile[13][21]~q ;
wire \rfile[12][21]~q ;
wire \Mux42~17_combout ;
wire \rfile[15][21]~q ;
wire \Mux42~18_combout ;
wire \rfile[9][21]~feeder_combout ;
wire \rfile[9][21]~q ;
wire \rfile[11][21]~feeder_combout ;
wire \rfile[11][21]~q ;
wire \rfile[8][21]~q ;
wire \rfile[10][21]~q ;
wire \Mux42~10_combout ;
wire \Mux42~11_combout ;
wire \rfile[7][21]~q ;
wire \rfile[6][21]~q ;
wire \rfile[5][21]~q ;
wire \Mux42~12_combout ;
wire \Mux42~13_combout ;
wire \rfile[2][21]~q ;
wire \rfile[3][21]~q ;
wire \rfile[1][21]~q ;
wire \Mux42~14_combout ;
wire \Mux42~15_combout ;
wire \Mux42~16_combout ;
wire \rfile[29][20]~q ;
wire \rfile[17][20]~q ;
wire \Mux43~0_combout ;
wire \rfile[21][20]~feeder_combout ;
wire \rfile[21][20]~q ;
wire \Mux43~1_combout ;
wire \rfile[28][20]~q ;
wire \rfile[16][20]~feeder_combout ;
wire \rfile[16][20]~q ;
wire \rfile[20][20]~feeder_combout ;
wire \rfile[20][20]~q ;
wire \Mux43~4_combout ;
wire \Mux43~5_combout ;
wire \rfile[30][20]~q ;
wire \rfile[26][20]~q ;
wire \rfile[18][20]~q ;
wire \Mux43~2_combout ;
wire \Mux43~3_combout ;
wire \Mux43~6_combout ;
wire \rfile[23][20]~q ;
wire \rfile[19][20]~q ;
wire \rfile[27][20]~q ;
wire \Mux43~7_combout ;
wire \rfile[31][20]~q ;
wire \Mux43~8_combout ;
wire \rfile[12][20]~q ;
wire \rfile[13][20]~feeder_combout ;
wire \rfile[13][20]~q ;
wire \Mux43~17_combout ;
wire \rfile[14][20]~q ;
wire \rfile[15][20]~q ;
wire \Mux43~18_combout ;
wire \rfile[2][20]~q ;
wire \rfile[3][20]~q ;
wire \Mux43~14_combout ;
wire \Mux43~15_combout ;
wire \rfile[9][20]~feeder_combout ;
wire \rfile[9][20]~q ;
wire \rfile[8][20]~q ;
wire \rfile[10][20]~q ;
wire \Mux43~12_combout ;
wire \Mux43~13_combout ;
wire \Mux43~16_combout ;
wire \rfile[7][20]~q ;
wire \rfile[4][20]~q ;
wire \rfile[5][20]~q ;
wire \Mux43~10_combout ;
wire \rfile[6][20]~feeder_combout ;
wire \rfile[6][20]~q ;
wire \Mux43~11_combout ;
wire \rfile[29][19]~q ;
wire \rfile[25][19]~q ;
wire \rfile[21][19]~q ;
wire \rfile[17][19]~q ;
wire \Mux44~0_combout ;
wire \Mux44~1_combout ;
wire \rfile[23][19]~q ;
wire \rfile[19][19]~q ;
wire \Mux44~7_combout ;
wire \rfile[31][19]~q ;
wire \rfile[27][19]~q ;
wire \Mux44~8_combout ;
wire \rfile[20][19]~q ;
wire \rfile[28][19]~q ;
wire \rfile[16][19]~q ;
wire \rfile[24][19]~q ;
wire \Mux44~4_combout ;
wire \Mux44~5_combout ;
wire \rfile[30][19]~q ;
wire \rfile[22][19]~q ;
wire \rfile[26][19]~q ;
wire \rfile[18][19]~feeder_combout ;
wire \rfile[18][19]~q ;
wire \Mux44~2_combout ;
wire \Mux44~3_combout ;
wire \Mux44~6_combout ;
wire \rfile[8][19]~q ;
wire \rfile[10][19]~q ;
wire \Mux44~10_combout ;
wire \rfile[11][19]~q ;
wire \rfile[9][19]~q ;
wire \Mux44~11_combout ;
wire \rfile[6][19]~q ;
wire \rfile[7][19]~q ;
wire \Mux44~13_combout ;
wire \rfile[1][19]~q ;
wire \rfile[3][19]~q ;
wire \Mux44~14_combout ;
wire \rfile[2][19]~q ;
wire \Mux44~15_combout ;
wire \Mux44~16_combout ;
wire \rfile[14][19]~feeder_combout ;
wire \rfile[14][19]~q ;
wire \rfile[15][19]~q ;
wire \rfile[13][19]~q ;
wire \rfile[12][19]~q ;
wire \Mux44~17_combout ;
wire \Mux44~18_combout ;
wire \rfile[21][18]~feeder_combout ;
wire \rfile[21][18]~q ;
wire \rfile[29][18]~q ;
wire \rfile[17][18]~q ;
wire \rfile[25][18]~q ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \rfile[23][18]~feeder_combout ;
wire \rfile[23][18]~q ;
wire \rfile[31][18]~q ;
wire \rfile[27][18]~q ;
wire \rfile[19][18]~feeder_combout ;
wire \rfile[19][18]~q ;
wire \Mux45~7_combout ;
wire \Mux45~8_combout ;
wire \rfile[30][18]~q ;
wire \rfile[26][18]~q ;
wire \rfile[18][18]~q ;
wire \rfile[22][18]~feeder_combout ;
wire \rfile[22][18]~q ;
wire \Mux45~2_combout ;
wire \Mux45~3_combout ;
wire \rfile[28][18]~q ;
wire \rfile[24][18]~q ;
wire \rfile[16][18]~q ;
wire \rfile[20][18]~q ;
wire \Mux45~4_combout ;
wire \Mux45~5_combout ;
wire \Mux45~6_combout ;
wire \rfile[4][18]~q ;
wire \Mux45~10_combout ;
wire \rfile[7][18]~q ;
wire \rfile[6][18]~feeder_combout ;
wire \rfile[6][18]~q ;
wire \Mux45~11_combout ;
wire \rfile[15][18]~q ;
wire \rfile[14][18]~q ;
wire \rfile[13][18]~q ;
wire \rfile[12][18]~q ;
wire \Mux45~17_combout ;
wire \Mux45~18_combout ;
wire \rfile[2][18]~q ;
wire \rfile[1][18]~q ;
wire \rfile[3][18]~feeder_combout ;
wire \rfile[3][18]~q ;
wire \Mux45~14_combout ;
wire \Mux45~15_combout ;
wire \rfile[11][18]~feeder_combout ;
wire \rfile[11][18]~q ;
wire \rfile[9][18]~q ;
wire \rfile[8][18]~q ;
wire \rfile[10][18]~feeder_combout ;
wire \rfile[10][18]~q ;
wire \Mux45~12_combout ;
wire \Mux45~13_combout ;
wire \Mux45~16_combout ;
wire \rfile[28][17]~q ;
wire \rfile[24][17]~q ;
wire \rfile[16][17]~q ;
wire \Mux46~4_combout ;
wire \Mux46~5_combout ;
wire \rfile[30][17]~q ;
wire \rfile[18][17]~q ;
wire \rfile[26][17]~q ;
wire \Mux46~2_combout ;
wire \Mux46~3_combout ;
wire \Mux46~6_combout ;
wire \rfile[27][17]~feeder_combout ;
wire \rfile[27][17]~q ;
wire \rfile[31][17]~q ;
wire \rfile[23][17]~q ;
wire \rfile[19][17]~feeder_combout ;
wire \rfile[19][17]~q ;
wire \Mux46~7_combout ;
wire \Mux46~8_combout ;
wire \rfile[29][17]~q ;
wire \rfile[25][17]~q ;
wire \rfile[17][17]~q ;
wire \rfile[21][17]~feeder_combout ;
wire \rfile[21][17]~q ;
wire \Mux46~0_combout ;
wire \Mux46~1_combout ;
wire \rfile[6][17]~feeder_combout ;
wire \rfile[6][17]~q ;
wire \rfile[7][17]~q ;
wire \rfile[5][17]~q ;
wire \rfile[4][17]~q ;
wire \Mux46~12_combout ;
wire \Mux46~13_combout ;
wire \rfile[3][17]~q ;
wire \rfile[1][17]~q ;
wire \Mux46~14_combout ;
wire \rfile[2][17]~feeder_combout ;
wire \rfile[2][17]~q ;
wire \Mux46~15_combout ;
wire \Mux46~16_combout ;
wire \rfile[9][17]~q ;
wire \rfile[11][17]~q ;
wire \rfile[10][17]~q ;
wire \rfile[8][17]~q ;
wire \Mux46~10_combout ;
wire \Mux46~11_combout ;
wire \rfile[15][17]~q ;
wire \rfile[14][17]~q ;
wire \rfile[12][17]~q ;
wire \rfile[13][17]~feeder_combout ;
wire \rfile[13][17]~q ;
wire \Mux46~17_combout ;
wire \Mux46~18_combout ;
wire \rfile[19][16]~q ;
wire \rfile[27][16]~q ;
wire \Mux47~7_combout ;
wire \rfile[23][16]~q ;
wire \rfile[31][16]~q ;
wire \Mux47~8_combout ;
wire \rfile[28][16]~q ;
wire \rfile[20][16]~feeder_combout ;
wire \rfile[20][16]~q ;
wire \rfile[16][16]~feeder_combout ;
wire \rfile[16][16]~q ;
wire \Mux47~4_combout ;
wire \Mux47~5_combout ;
wire \rfile[30][16]~q ;
wire \rfile[26][16]~q ;
wire \Mux47~3_combout ;
wire \Mux47~6_combout ;
wire \rfile[29][16]~q ;
wire \rfile[21][16]~feeder_combout ;
wire \rfile[21][16]~q ;
wire \rfile[17][16]~q ;
wire \rfile[25][16]~q ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \rfile[9][16]~feeder_combout ;
wire \rfile[9][16]~q ;
wire \rfile[11][16]~q ;
wire \rfile[10][16]~q ;
wire \Mux47~12_combout ;
wire \Mux47~13_combout ;
wire \rfile[1][16]~q ;
wire \rfile[3][16]~q ;
wire \Mux47~14_combout ;
wire \rfile[2][16]~feeder_combout ;
wire \rfile[2][16]~q ;
wire \Mux47~15_combout ;
wire \Mux47~16_combout ;
wire \rfile[6][16]~feeder_combout ;
wire \rfile[6][16]~q ;
wire \rfile[7][16]~q ;
wire \rfile[5][16]~q ;
wire \Mux47~10_combout ;
wire \Mux47~11_combout ;
wire \rfile[14][16]~feeder_combout ;
wire \rfile[14][16]~q ;
wire \rfile[15][16]~feeder_combout ;
wire \rfile[15][16]~q ;
wire \rfile[12][16]~q ;
wire \rfile[13][16]~feeder_combout ;
wire \rfile[13][16]~q ;
wire \Mux47~17_combout ;
wire \Mux47~18_combout ;
wire \rfile[21][15]~q ;
wire \rfile[17][15]~feeder_combout ;
wire \rfile[17][15]~q ;
wire \Mux48~0_combout ;
wire \rfile[25][15]~q ;
wire \rfile[29][15]~q ;
wire \Mux48~1_combout ;
wire \rfile[27][15]~q ;
wire \rfile[31][15]~q ;
wire \rfile[23][15]~q ;
wire \rfile[19][15]~q ;
wire \Mux48~7_combout ;
wire \Mux48~8_combout ;
wire \rfile[30][15]~feeder_combout ;
wire \rfile[30][15]~q ;
wire \rfile[22][15]~q ;
wire \rfile[18][15]~q ;
wire \rfile[26][15]~q ;
wire \Mux48~2_combout ;
wire \Mux48~3_combout ;
wire \rfile[20][15]~q ;
wire \rfile[16][15]~q ;
wire \Mux48~4_combout ;
wire \Mux48~5_combout ;
wire \Mux48~6_combout ;
wire \rfile[14][15]~feeder_combout ;
wire \rfile[14][15]~q ;
wire \rfile[15][15]~feeder_combout ;
wire \rfile[15][15]~q ;
wire \rfile[12][15]~q ;
wire \rfile[13][15]~q ;
wire \Mux48~17_combout ;
wire \Mux48~18_combout ;
wire \rfile[9][15]~q ;
wire \rfile[11][15]~q ;
wire \rfile[10][15]~q ;
wire \rfile[8][15]~q ;
wire \Mux48~10_combout ;
wire \Mux48~11_combout ;
wire \rfile[2][15]~feeder_combout ;
wire \rfile[2][15]~q ;
wire \rfile[3][15]~q ;
wire \rfile[1][15]~q ;
wire \Mux48~14_combout ;
wire \Mux48~15_combout ;
wire \rfile[7][15]~q ;
wire \rfile[6][15]~q ;
wire \rfile[5][15]~feeder_combout ;
wire \rfile[5][15]~q ;
wire \rfile[4][15]~feeder_combout ;
wire \rfile[4][15]~q ;
wire \Mux48~12_combout ;
wire \Mux48~13_combout ;
wire \Mux48~16_combout ;
wire \rfile[31][14]~q ;
wire \rfile[23][14]~q ;
wire \rfile[27][14]~q ;
wire \rfile[19][14]~q ;
wire \Mux49~7_combout ;
wire \Mux49~8_combout ;
wire \rfile[30][14]~q ;
wire \rfile[26][14]~q ;
wire \rfile[18][14]~q ;
wire \rfile[22][14]~q ;
wire \Mux49~2_combout ;
wire \Mux49~3_combout ;
wire \rfile[28][14]~q ;
wire \rfile[20][14]~q ;
wire \rfile[16][14]~q ;
wire \Mux49~4_combout ;
wire \Mux49~5_combout ;
wire \Mux49~6_combout ;
wire \rfile[21][14]~feeder_combout ;
wire \rfile[21][14]~q ;
wire \rfile[29][14]~feeder_combout ;
wire \rfile[29][14]~q ;
wire \rfile[17][14]~q ;
wire \rfile[25][14]~feeder_combout ;
wire \rfile[25][14]~q ;
wire \Mux49~0_combout ;
wire \Mux49~1_combout ;
wire \rfile[14][14]~feeder_combout ;
wire \rfile[14][14]~q ;
wire \rfile[15][14]~feeder_combout ;
wire \rfile[15][14]~q ;
wire \rfile[12][14]~q ;
wire \rfile[13][14]~feeder_combout ;
wire \rfile[13][14]~q ;
wire \Mux49~17_combout ;
wire \Mux49~18_combout ;
wire \rfile[2][14]~feeder_combout ;
wire \rfile[2][14]~q ;
wire \rfile[1][14]~q ;
wire \rfile[3][14]~q ;
wire \Mux49~14_combout ;
wire \Mux49~15_combout ;
wire \rfile[11][14]~feeder_combout ;
wire \rfile[11][14]~q ;
wire \rfile[9][14]~q ;
wire \rfile[10][14]~q ;
wire \rfile[8][14]~q ;
wire \Mux49~12_combout ;
wire \Mux49~13_combout ;
wire \Mux49~16_combout ;
wire \rfile[7][14]~feeder_combout ;
wire \rfile[7][14]~q ;
wire \rfile[6][14]~feeder_combout ;
wire \rfile[6][14]~q ;
wire \rfile[4][14]~q ;
wire \rfile[5][14]~feeder_combout ;
wire \rfile[5][14]~q ;
wire \Mux49~10_combout ;
wire \Mux49~11_combout ;
wire \rfile[30][13]~q ;
wire \rfile[22][13]~q ;
wire \rfile[18][13]~q ;
wire \rfile[26][13]~q ;
wire \Mux50~2_combout ;
wire \Mux50~3_combout ;
wire \rfile[28][13]~q ;
wire \rfile[16][13]~q ;
wire \rfile[24][13]~q ;
wire \Mux50~4_combout ;
wire \Mux50~5_combout ;
wire \Mux50~6_combout ;
wire \rfile[25][13]~feeder_combout ;
wire \rfile[25][13]~q ;
wire \rfile[29][13]~q ;
wire \rfile[21][13]~q ;
wire \rfile[17][13]~q ;
wire \Mux50~0_combout ;
wire \Mux50~1_combout ;
wire \rfile[27][13]~feeder_combout ;
wire \rfile[27][13]~q ;
wire \rfile[31][13]~q ;
wire \rfile[23][13]~q ;
wire \rfile[19][13]~q ;
wire \Mux50~7_combout ;
wire \Mux50~8_combout ;
wire \rfile[1][13]~q ;
wire \rfile[3][13]~feeder_combout ;
wire \rfile[3][13]~q ;
wire \Mux50~14_combout ;
wire \rfile[2][13]~q ;
wire \Mux50~15_combout ;
wire \rfile[6][13]~q ;
wire \rfile[4][13]~q ;
wire \rfile[5][13]~q ;
wire \Mux50~12_combout ;
wire \Mux50~13_combout ;
wire \Mux50~16_combout ;
wire \rfile[11][13]~q ;
wire \rfile[9][13]~q ;
wire \rfile[8][13]~q ;
wire \rfile[10][13]~q ;
wire \Mux50~10_combout ;
wire \Mux50~11_combout ;
wire \rfile[15][13]~feeder_combout ;
wire \rfile[15][13]~q ;
wire \rfile[14][13]~feeder_combout ;
wire \rfile[14][13]~q ;
wire \rfile[13][13]~q ;
wire \rfile[12][13]~q ;
wire \Mux50~17_combout ;
wire \Mux50~18_combout ;
wire \rfile[31][12]~q ;
wire \rfile[19][12]~q ;
wire \rfile[27][12]~q ;
wire \Mux51~7_combout ;
wire \rfile[23][12]~q ;
wire \Mux51~8_combout ;
wire \rfile[21][12]~feeder_combout ;
wire \rfile[21][12]~q ;
wire \rfile[29][12]~q ;
wire \rfile[17][12]~q ;
wire \rfile[25][12]~q ;
wire \Mux51~0_combout ;
wire \Mux51~1_combout ;
wire \rfile[28][12]~q ;
wire \rfile[20][12]~feeder_combout ;
wire \rfile[20][12]~q ;
wire \rfile[16][12]~feeder_combout ;
wire \rfile[16][12]~q ;
wire \Mux51~4_combout ;
wire \Mux51~5_combout ;
wire \rfile[26][12]~q ;
wire \rfile[22][12]~q ;
wire \rfile[18][12]~q ;
wire \Mux51~2_combout ;
wire \Mux51~3_combout ;
wire \Mux51~6_combout ;
wire \rfile[15][12]~feeder_combout ;
wire \rfile[15][12]~q ;
wire \rfile[14][12]~q ;
wire \rfile[13][12]~q ;
wire \rfile[12][12]~q ;
wire \Mux51~17_combout ;
wire \Mux51~18_combout ;
wire \rfile[5][12]~q ;
wire \Mux51~10_combout ;
wire \rfile[6][12]~q ;
wire \rfile[7][12]~q ;
wire \Mux51~11_combout ;
wire \rfile[2][12]~q ;
wire \rfile[3][12]~q ;
wire \rfile[1][12]~q ;
wire \Mux51~14_combout ;
wire \Mux51~15_combout ;
wire \rfile[11][12]~q ;
wire \rfile[9][12]~feeder_combout ;
wire \rfile[9][12]~q ;
wire \Mux51~13_combout ;
wire \Mux51~16_combout ;
wire \rfile[17][9]~q ;
wire \rfile[21][9]~q ;
wire \Mux54~0_combout ;
wire \rfile[29][9]~q ;
wire \rfile[25][9]~q ;
wire \Mux54~1_combout ;
wire \rfile[27][9]~feeder_combout ;
wire \rfile[27][9]~q ;
wire \rfile[31][9]~q ;
wire \rfile[23][9]~feeder_combout ;
wire \rfile[23][9]~q ;
wire \rfile[19][9]~q ;
wire \Mux54~7_combout ;
wire \Mux54~8_combout ;
wire \rfile[30][9]~q ;
wire \rfile[22][9]~q ;
wire \rfile[26][9]~q ;
wire \rfile[18][9]~q ;
wire \Mux54~2_combout ;
wire \Mux54~3_combout ;
wire \rfile[28][9]~q ;
wire \rfile[16][9]~q ;
wire \rfile[24][9]~q ;
wire \Mux54~4_combout ;
wire \Mux54~5_combout ;
wire \Mux54~6_combout ;
wire \rfile[15][9]~feeder_combout ;
wire \rfile[15][9]~q ;
wire \rfile[14][9]~feeder_combout ;
wire \rfile[14][9]~q ;
wire \rfile[12][9]~q ;
wire \rfile[13][9]~q ;
wire \Mux54~17_combout ;
wire \Mux54~18_combout ;
wire \rfile[11][9]~q ;
wire \rfile[9][9]~q ;
wire \rfile[8][9]~q ;
wire \rfile[10][9]~q ;
wire \Mux54~10_combout ;
wire \Mux54~11_combout ;
wire \rfile[1][9]~q ;
wire \rfile[3][9]~q ;
wire \Mux54~14_combout ;
wire \Mux54~15_combout ;
wire \rfile[6][9]~q ;
wire \rfile[7][9]~q ;
wire \Mux54~13_combout ;
wire \Mux54~16_combout ;
wire \rfile[31][8]~q ;
wire \rfile[23][8]~q ;
wire \rfile[19][8]~q ;
wire \rfile[27][8]~q ;
wire \Mux55~7_combout ;
wire \Mux55~8_combout ;
wire \rfile[26][8]~q ;
wire \rfile[18][8]~q ;
wire \rfile[22][8]~q ;
wire \Mux55~2_combout ;
wire \Mux55~3_combout ;
wire \rfile[24][8]~q ;
wire \rfile[16][8]~feeder_combout ;
wire \rfile[16][8]~q ;
wire \rfile[20][8]~feeder_combout ;
wire \rfile[20][8]~q ;
wire \Mux55~4_combout ;
wire \Mux55~5_combout ;
wire \Mux55~6_combout ;
wire \rfile[29][8]~q ;
wire \rfile[21][8]~feeder_combout ;
wire \rfile[21][8]~q ;
wire \rfile[25][8]~q ;
wire \rfile[17][8]~q ;
wire \Mux55~0_combout ;
wire \Mux55~1_combout ;
wire \rfile[15][8]~q ;
wire \rfile[14][8]~feeder_combout ;
wire \rfile[14][8]~q ;
wire \rfile[12][8]~q ;
wire \rfile[13][8]~q ;
wire \Mux55~17_combout ;
wire \Mux55~18_combout ;
wire \rfile[6][8]~feeder_combout ;
wire \rfile[6][8]~q ;
wire \rfile[5][8]~q ;
wire \rfile[4][8]~q ;
wire \Mux55~10_combout ;
wire \rfile[7][8]~feeder_combout ;
wire \rfile[7][8]~q ;
wire \Mux55~11_combout ;
wire \rfile[11][8]~q ;
wire \rfile[9][8]~q ;
wire \rfile[8][8]~q ;
wire \rfile[10][8]~q ;
wire \Mux55~12_combout ;
wire \Mux55~13_combout ;
wire \rfile[2][8]~feeder_combout ;
wire \rfile[2][8]~q ;
wire \rfile[3][8]~q ;
wire \rfile[1][8]~q ;
wire \Mux55~14_combout ;
wire \Mux55~15_combout ;
wire \Mux55~16_combout ;
wire \rfile[27][11]~feeder_combout ;
wire \rfile[27][11]~q ;
wire \rfile[31][11]~q ;
wire \rfile[23][11]~feeder_combout ;
wire \rfile[23][11]~q ;
wire \rfile[19][11]~feeder_combout ;
wire \rfile[19][11]~q ;
wire \Mux52~7_combout ;
wire \Mux52~8_combout ;
wire \rfile[29][11]~feeder_combout ;
wire \rfile[29][11]~q ;
wire \rfile[17][11]~q ;
wire \rfile[21][11]~q ;
wire \Mux52~0_combout ;
wire \rfile[25][11]~feeder_combout ;
wire \rfile[25][11]~q ;
wire \Mux52~1_combout ;
wire \rfile[18][11]~feeder_combout ;
wire \rfile[18][11]~q ;
wire \Mux52~2_combout ;
wire \rfile[22][11]~feeder_combout ;
wire \rfile[22][11]~q ;
wire \Mux52~3_combout ;
wire \rfile[20][11]~feeder_combout ;
wire \rfile[20][11]~q ;
wire \rfile[24][11]~q ;
wire \rfile[16][11]~q ;
wire \Mux52~4_combout ;
wire \rfile[28][11]~q ;
wire \Mux52~5_combout ;
wire \Mux52~6_combout ;
wire \rfile[15][11]~q ;
wire \rfile[14][11]~feeder_combout ;
wire \rfile[14][11]~q ;
wire \rfile[12][11]~q ;
wire \rfile[13][11]~feeder_combout ;
wire \rfile[13][11]~q ;
wire \Mux52~17_combout ;
wire \Mux52~18_combout ;
wire \rfile[7][11]~q ;
wire \rfile[4][11]~q ;
wire \rfile[5][11]~q ;
wire \Mux52~12_combout ;
wire \Mux52~13_combout ;
wire \rfile[2][11]~q ;
wire \rfile[1][11]~q ;
wire \rfile[3][11]~feeder_combout ;
wire \rfile[3][11]~q ;
wire \Mux52~14_combout ;
wire \Mux52~15_combout ;
wire \Mux52~16_combout ;
wire \rfile[9][11]~feeder_combout ;
wire \rfile[9][11]~q ;
wire \rfile[11][11]~q ;
wire \rfile[10][11]~q ;
wire \rfile[8][11]~q ;
wire \Mux52~10_combout ;
wire \Mux52~11_combout ;
wire \rfile[25][10]~q ;
wire \Mux53~0_combout ;
wire \rfile[21][10]~q ;
wire \rfile[29][10]~feeder_combout ;
wire \rfile[29][10]~q ;
wire \Mux53~1_combout ;
wire \rfile[23][10]~feeder_combout ;
wire \rfile[23][10]~q ;
wire \rfile[31][10]~q ;
wire \rfile[27][10]~feeder_combout ;
wire \rfile[27][10]~q ;
wire \rfile[19][10]~feeder_combout ;
wire \rfile[19][10]~q ;
wire \Mux53~7_combout ;
wire \Mux53~8_combout ;
wire \rfile[28][10]~q ;
wire \rfile[24][10]~feeder_combout ;
wire \rfile[24][10]~q ;
wire \rfile[20][10]~q ;
wire \rfile[16][10]~q ;
wire \Mux53~4_combout ;
wire \Mux53~5_combout ;
wire \rfile[30][10]~q ;
wire \rfile[18][10]~feeder_combout ;
wire \rfile[18][10]~q ;
wire \rfile[22][10]~feeder_combout ;
wire \rfile[22][10]~q ;
wire \Mux53~2_combout ;
wire \Mux53~3_combout ;
wire \Mux53~6_combout ;
wire \rfile[6][10]~q ;
wire \rfile[7][10]~q ;
wire \rfile[4][10]~q ;
wire \rfile[5][10]~q ;
wire \Mux53~10_combout ;
wire \Mux53~11_combout ;
wire \rfile[15][10]~q ;
wire \rfile[14][10]~feeder_combout ;
wire \rfile[14][10]~q ;
wire \rfile[13][10]~feeder_combout ;
wire \rfile[13][10]~q ;
wire \rfile[12][10]~q ;
wire \Mux53~17_combout ;
wire \Mux53~18_combout ;
wire \rfile[11][10]~feeder_combout ;
wire \rfile[11][10]~q ;
wire \rfile[9][10]~feeder_combout ;
wire \rfile[9][10]~q ;
wire \rfile[8][10]~q ;
wire \rfile[10][10]~q ;
wire \Mux53~12_combout ;
wire \Mux53~13_combout ;
wire \rfile[2][10]~feeder_combout ;
wire \rfile[2][10]~q ;
wire \rfile[3][10]~feeder_combout ;
wire \rfile[3][10]~q ;
wire \rfile[1][10]~feeder_combout ;
wire \rfile[1][10]~q ;
wire \Mux53~14_combout ;
wire \Mux53~15_combout ;
wire \Mux53~16_combout ;
wire \rfile[17][7]~feeder_combout ;
wire \rfile[17][7]~q ;
wire \rfile[21][7]~q ;
wire \Mux56~0_combout ;
wire \rfile[29][7]~q ;
wire \rfile[25][7]~q ;
wire \Mux56~1_combout ;
wire \rfile[31][7]~q ;
wire \rfile[27][7]~q ;
wire \rfile[19][7]~q ;
wire \rfile[23][7]~q ;
wire \Mux56~7_combout ;
wire \Mux56~8_combout ;
wire \rfile[28][7]~feeder_combout ;
wire \rfile[28][7]~q ;
wire \rfile[20][7]~q ;
wire \rfile[24][7]~feeder_combout ;
wire \rfile[24][7]~q ;
wire \rfile[16][7]~feeder_combout ;
wire \rfile[16][7]~q ;
wire \Mux56~4_combout ;
wire \Mux56~5_combout ;
wire \rfile[22][7]~q ;
wire \rfile[30][7]~q ;
wire \rfile[26][7]~feeder_combout ;
wire \rfile[26][7]~q ;
wire \rfile[18][7]~feeder_combout ;
wire \rfile[18][7]~q ;
wire \Mux56~2_combout ;
wire \Mux56~3_combout ;
wire \Mux56~6_combout ;
wire \rfile[15][7]~feeder_combout ;
wire \rfile[15][7]~q ;
wire \rfile[14][7]~q ;
wire \rfile[13][7]~q ;
wire \Mux56~17_combout ;
wire \Mux56~18_combout ;
wire \rfile[4][7]~q ;
wire \rfile[5][7]~q ;
wire \Mux56~12_combout ;
wire \rfile[7][7]~q ;
wire \Mux56~13_combout ;
wire \rfile[3][7]~q ;
wire \rfile[1][7]~q ;
wire \Mux56~14_combout ;
wire \Mux56~15_combout ;
wire \Mux56~16_combout ;
wire \rfile[10][7]~q ;
wire \rfile[8][7]~q ;
wire \Mux56~10_combout ;
wire \rfile[11][7]~q ;
wire \rfile[9][7]~feeder_combout ;
wire \rfile[9][7]~q ;
wire \Mux56~11_combout ;
wire \rfile[21][6]~feeder_combout ;
wire \rfile[21][6]~q ;
wire \rfile[29][6]~feeder_combout ;
wire \rfile[29][6]~q ;
wire \rfile[25][6]~q ;
wire \rfile[17][6]~q ;
wire \Mux57~0_combout ;
wire \Mux57~1_combout ;
wire \rfile[24][6]~q ;
wire \rfile[20][6]~q ;
wire \rfile[16][6]~q ;
wire \Mux57~4_combout ;
wire \rfile[28][6]~feeder_combout ;
wire \rfile[28][6]~q ;
wire \Mux57~5_combout ;
wire \rfile[30][6]~q ;
wire \rfile[22][6]~feeder_combout ;
wire \rfile[22][6]~q ;
wire \rfile[18][6]~q ;
wire \Mux57~2_combout ;
wire \Mux57~3_combout ;
wire \Mux57~6_combout ;
wire \rfile[31][6]~feeder_combout ;
wire \rfile[31][6]~q ;
wire \rfile[23][6]~q ;
wire \rfile[27][6]~q ;
wire \rfile[19][6]~q ;
wire \Mux57~7_combout ;
wire \Mux57~8_combout ;
wire \rfile[7][6]~feeder_combout ;
wire \rfile[7][6]~q ;
wire \rfile[5][6]~q ;
wire \Mux57~10_combout ;
wire \rfile[6][6]~feeder_combout ;
wire \rfile[6][6]~q ;
wire \Mux57~11_combout ;
wire \rfile[14][6]~feeder_combout ;
wire \rfile[14][6]~q ;
wire \rfile[12][6]~q ;
wire \rfile[13][6]~q ;
wire \Mux57~17_combout ;
wire \rfile[15][6]~feeder_combout ;
wire \rfile[15][6]~q ;
wire \Mux57~18_combout ;
wire \rfile[2][6]~feeder_combout ;
wire \rfile[2][6]~q ;
wire \rfile[1][6]~feeder_combout ;
wire \rfile[1][6]~q ;
wire \rfile[3][6]~feeder_combout ;
wire \rfile[3][6]~q ;
wire \Mux57~14_combout ;
wire \Mux57~15_combout ;
wire \rfile[9][6]~q ;
wire \rfile[10][6]~q ;
wire \rfile[8][6]~q ;
wire \Mux57~12_combout ;
wire \Mux57~13_combout ;
wire \Mux57~16_combout ;
wire \rfile[27][5]~feeder_combout ;
wire \rfile[27][5]~q ;
wire \rfile[19][5]~feeder_combout ;
wire \rfile[19][5]~q ;
wire \rfile[23][5]~feeder_combout ;
wire \rfile[23][5]~q ;
wire \Mux58~7_combout ;
wire \rfile[31][5]~feeder_combout ;
wire \rfile[31][5]~q ;
wire \Mux58~8_combout ;
wire \rfile[17][5]~q ;
wire \rfile[21][5]~q ;
wire \Mux58~0_combout ;
wire \rfile[29][5]~q ;
wire \rfile[25][5]~q ;
wire \Mux58~1_combout ;
wire \rfile[20][5]~q ;
wire \rfile[24][5]~q ;
wire \rfile[16][5]~q ;
wire \Mux58~4_combout ;
wire \Mux58~5_combout ;
wire \rfile[30][5]~q ;
wire \rfile[26][5]~q ;
wire \Mux58~2_combout ;
wire \Mux58~3_combout ;
wire \Mux58~6_combout ;
wire \rfile[11][5]~feeder_combout ;
wire \rfile[11][5]~q ;
wire \rfile[10][5]~q ;
wire \rfile[8][5]~q ;
wire \Mux58~10_combout ;
wire \rfile[9][5]~feeder_combout ;
wire \rfile[9][5]~q ;
wire \Mux58~11_combout ;
wire \rfile[15][5]~feeder_combout ;
wire \rfile[15][5]~q ;
wire \rfile[14][5]~q ;
wire \rfile[13][5]~q ;
wire \rfile[12][5]~q ;
wire \Mux58~17_combout ;
wire \Mux58~18_combout ;
wire \rfile[3][5]~feeder_combout ;
wire \rfile[3][5]~q ;
wire \rfile[1][5]~feeder_combout ;
wire \rfile[1][5]~q ;
wire \Mux58~14_combout ;
wire \rfile[2][5]~feeder_combout ;
wire \rfile[2][5]~q ;
wire \Mux58~15_combout ;
wire \rfile[6][5]~feeder_combout ;
wire \rfile[6][5]~q ;
wire \rfile[7][5]~feeder_combout ;
wire \rfile[7][5]~q ;
wire \rfile[5][5]~q ;
wire \rfile[4][5]~q ;
wire \Mux58~12_combout ;
wire \Mux58~13_combout ;
wire \Mux58~16_combout ;
wire \rfile[21][2]~q ;
wire \rfile[17][2]~feeder_combout ;
wire \rfile[17][2]~q ;
wire \Mux29~0_combout ;
wire \rfile[29][2]~q ;
wire \rfile[25][2]~q ;
wire \Mux29~1_combout ;
wire \rfile[23][2]~feeder_combout ;
wire \rfile[23][2]~q ;
wire \rfile[19][2]~q ;
wire \Mux29~7_combout ;
wire \rfile[31][2]~q ;
wire \rfile[27][2]~q ;
wire \Mux29~8_combout ;
wire \rfile[30][2]~q ;
wire \rfile[22][2]~feeder_combout ;
wire \rfile[22][2]~q ;
wire \rfile[18][2]~feeder_combout ;
wire \rfile[18][2]~q ;
wire \rfile[26][2]~feeder_combout ;
wire \rfile[26][2]~q ;
wire \Mux29~2_combout ;
wire \Mux29~3_combout ;
wire \rfile[20][2]~q ;
wire \rfile[16][2]~feeder_combout ;
wire \rfile[16][2]~q ;
wire \rfile[24][2]~feeder_combout ;
wire \rfile[24][2]~q ;
wire \Mux29~4_combout ;
wire \Mux29~5_combout ;
wire \Mux29~6_combout ;
wire \rfile[9][2]~feeder_combout ;
wire \rfile[9][2]~q ;
wire \rfile[11][2]~feeder_combout ;
wire \rfile[11][2]~q ;
wire \rfile[10][2]~q ;
wire \rfile[8][2]~feeder_combout ;
wire \rfile[8][2]~q ;
wire \Mux29~10_combout ;
wire \Mux29~11_combout ;
wire \rfile[15][2]~feeder_combout ;
wire \rfile[15][2]~q ;
wire \rfile[14][2]~q ;
wire \rfile[13][2]~feeder_combout ;
wire \rfile[13][2]~q ;
wire \rfile[12][2]~q ;
wire \Mux29~17_combout ;
wire \Mux29~18_combout ;
wire \rfile[6][2]~q ;
wire \rfile[7][2]~q ;
wire \rfile[5][2]~q ;
wire \rfile[4][2]~q ;
wire \Mux29~12_combout ;
wire \Mux29~13_combout ;
wire \rfile[2][2]~feeder_combout ;
wire \rfile[2][2]~q ;
wire \rfile[1][2]~q ;
wire \rfile[3][2]~feeder_combout ;
wire \rfile[3][2]~q ;
wire \Mux29~14_combout ;
wire \Mux29~15_combout ;
wire \Mux29~16_combout ;
wire \rfile[16][1]~q ;
wire \rfile[24][1]~q ;
wire \Mux30~4_combout ;
wire \rfile[20][1]~q ;
wire \rfile[28][1]~feeder_combout ;
wire \rfile[28][1]~q ;
wire \Mux30~5_combout ;
wire \rfile[22][1]~q ;
wire \rfile[30][1]~q ;
wire \Mux30~3_combout ;
wire \Mux30~6_combout ;
wire \rfile[27][1]~q ;
wire \rfile[31][1]~q ;
wire \rfile[23][1]~feeder_combout ;
wire \rfile[23][1]~q ;
wire \rfile[19][1]~feeder_combout ;
wire \rfile[19][1]~q ;
wire \Mux30~7_combout ;
wire \Mux30~8_combout ;
wire \rfile[25][1]~q ;
wire \rfile[29][1]~q ;
wire \rfile[17][1]~q ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \rfile[11][1]~q ;
wire \rfile[9][1]~q ;
wire \rfile[10][1]~q ;
wire \rfile[8][1]~q ;
wire \Mux30~10_combout ;
wire \Mux30~11_combout ;
wire \rfile[15][1]~q ;
wire \rfile[14][1]~q ;
wire \rfile[13][1]~feeder_combout ;
wire \rfile[13][1]~q ;
wire \Mux30~17_combout ;
wire \Mux30~18_combout ;
wire \rfile[7][1]~feeder_combout ;
wire \rfile[7][1]~q ;
wire \rfile[6][1]~q ;
wire \Mux30~13_combout ;
wire \rfile[1][1]~q ;
wire \rfile[3][1]~q ;
wire \Mux30~14_combout ;
wire \Mux30~15_combout ;
wire \Mux30~16_combout ;
wire \rfile[29][0]~q ;
wire \rfile[21][0]~q ;
wire \rfile[25][0]~q ;
wire \rfile[17][0]~q ;
wire \Mux63~0_combout ;
wire \Mux63~1_combout ;
wire \rfile[23][0]~q ;
wire \rfile[31][0]~q ;
wire \rfile[27][0]~q ;
wire \rfile[19][0]~q ;
wire \Mux63~7_combout ;
wire \Mux63~8_combout ;
wire \rfile[18][0]~q ;
wire \rfile[22][0]~q ;
wire \Mux63~2_combout ;
wire \rfile[30][0]~q ;
wire \rfile[26][0]~q ;
wire \Mux63~3_combout ;
wire \rfile[24][0]~q ;
wire \rfile[20][0]~q ;
wire \rfile[16][0]~q ;
wire \Mux63~4_combout ;
wire \Mux63~5_combout ;
wire \Mux63~6_combout ;
wire \rfile[3][0]~q ;
wire \rfile[1][0]~q ;
wire \Mux63~14_combout ;
wire \rfile[2][0]~feeder_combout ;
wire \rfile[2][0]~q ;
wire \Mux63~15_combout ;
wire \rfile[11][0]~q ;
wire \rfile[9][0]~q ;
wire \rfile[10][0]~q ;
wire \rfile[8][0]~q ;
wire \Mux63~12_combout ;
wire \Mux63~13_combout ;
wire \Mux63~16_combout ;
wire \rfile[13][0]~q ;
wire \Mux63~17_combout ;
wire \rfile[14][0]~q ;
wire \rfile[15][0]~q ;
wire \Mux63~18_combout ;
wire \rfile[7][0]~q ;
wire \rfile[6][0]~q ;
wire \rfile[5][0]~q ;
wire \rfile[4][0]~q ;
wire \Mux63~10_combout ;
wire \Mux63~11_combout ;
wire \rfile[21][1]~q ;
wire \Mux62~0_combout ;
wire \Mux62~1_combout ;
wire \Mux62~4_combout ;
wire \Mux62~5_combout ;
wire \Mux62~3_combout ;
wire \Mux62~6_combout ;
wire \Mux62~7_combout ;
wire \Mux62~8_combout ;
wire \Mux62~10_combout ;
wire \Mux62~11_combout ;
wire \Mux62~17_combout ;
wire \Mux62~18_combout ;
wire \Mux62~14_combout ;
wire \Mux62~15_combout ;
wire \rfile[5][1]~q ;
wire \Mux62~12_combout ;
wire \Mux62~13_combout ;
wire \Mux62~16_combout ;
wire \rfile[23][4]~q ;
wire \rfile[31][4]~q ;
wire \rfile[27][4]~q ;
wire \rfile[19][4]~q ;
wire \Mux27~7_combout ;
wire \Mux27~8_combout ;
wire \rfile[25][4]~q ;
wire \rfile[17][4]~feeder_combout ;
wire \rfile[17][4]~q ;
wire \Mux27~0_combout ;
wire \rfile[21][4]~q ;
wire \rfile[29][4]~q ;
wire \Mux27~1_combout ;
wire \rfile[26][4]~feeder_combout ;
wire \rfile[26][4]~q ;
wire \rfile[22][4]~feeder_combout ;
wire \rfile[22][4]~q ;
wire \rfile[18][4]~q ;
wire \Mux27~2_combout ;
wire \Mux27~3_combout ;
wire \rfile[24][4]~q ;
wire \rfile[28][4]~q ;
wire \rfile[20][4]~q ;
wire \rfile[16][4]~feeder_combout ;
wire \rfile[16][4]~q ;
wire \Mux27~4_combout ;
wire \Mux27~5_combout ;
wire \Mux27~6_combout ;
wire \rfile[15][4]~q ;
wire \rfile[14][4]~q ;
wire \rfile[13][4]~q ;
wire \rfile[12][4]~q ;
wire \Mux27~17_combout ;
wire \Mux27~18_combout ;
wire \rfile[7][4]~q ;
wire \rfile[6][4]~q ;
wire \rfile[5][4]~q ;
wire \rfile[4][4]~q ;
wire \Mux27~10_combout ;
wire \Mux27~11_combout ;
wire \rfile[3][4]~q ;
wire \rfile[1][4]~q ;
wire \Mux27~14_combout ;
wire \rfile[2][4]~feeder_combout ;
wire \rfile[2][4]~q ;
wire \Mux27~15_combout ;
wire \rfile[11][4]~feeder_combout ;
wire \rfile[11][4]~q ;
wire \rfile[9][4]~q ;
wire \rfile[10][4]~q ;
wire \rfile[8][4]~q ;
wire \Mux27~12_combout ;
wire \Mux27~13_combout ;
wire \Mux27~16_combout ;
wire \rfile[23][3]~feeder_combout ;
wire \rfile[23][3]~q ;
wire \rfile[31][3]~q ;
wire \rfile[27][3]~q ;
wire \Mux28~7_combout ;
wire \Mux28~8_combout ;
wire \rfile[21][3]~feeder_combout ;
wire \rfile[21][3]~q ;
wire \rfile[29][3]~feeder_combout ;
wire \rfile[29][3]~q ;
wire \rfile[25][3]~q ;
wire \rfile[17][3]~feeder_combout ;
wire \rfile[17][3]~q ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \rfile[30][3]~q ;
wire \rfile[22][3]~q ;
wire \rfile[18][3]~feeder_combout ;
wire \rfile[18][3]~q ;
wire \Mux28~2_combout ;
wire \rfile[26][3]~q ;
wire \Mux28~3_combout ;
wire \rfile[16][3]~q ;
wire \rfile[20][3]~feeder_combout ;
wire \rfile[20][3]~q ;
wire \Mux28~4_combout ;
wire \rfile[24][3]~q ;
wire \Mux28~5_combout ;
wire \Mux28~6_combout ;
wire \rfile[14][3]~q ;
wire \rfile[12][3]~q ;
wire \rfile[13][3]~q ;
wire \Mux28~17_combout ;
wire \rfile[15][3]~feeder_combout ;
wire \rfile[15][3]~q ;
wire \Mux28~18_combout ;
wire \rfile[7][3]~q ;
wire \rfile[4][3]~q ;
wire \rfile[5][3]~q ;
wire \Mux28~10_combout ;
wire \rfile[6][3]~q ;
wire \Mux28~11_combout ;
wire \rfile[3][3]~q ;
wire \rfile[1][3]~feeder_combout ;
wire \rfile[1][3]~q ;
wire \Mux28~14_combout ;
wire \rfile[2][3]~q ;
wire \Mux28~15_combout ;
wire \rfile[11][3]~q ;
wire \rfile[9][3]~feeder_combout ;
wire \rfile[9][3]~q ;
wire \rfile[10][3]~q ;
wire \Mux28~12_combout ;
wire \Mux28~13_combout ;
wire \Mux28~16_combout ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \Mux61~7_combout ;
wire \Mux61~8_combout ;
wire \Mux61~4_combout ;
wire \rfile[28][2]~feeder_combout ;
wire \rfile[28][2]~q ;
wire \Mux61~5_combout ;
wire \Mux61~2_combout ;
wire \Mux61~3_combout ;
wire \Mux61~6_combout ;
wire \Mux61~12_combout ;
wire \Mux61~13_combout ;
wire \Mux61~14_combout ;
wire \Mux61~15_combout ;
wire \Mux61~16_combout ;
wire \Mux61~10_combout ;
wire \Mux61~11_combout ;
wire \Mux61~17_combout ;
wire \Mux61~18_combout ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \Mux23~7_combout ;
wire \Mux23~8_combout ;
wire \rfile[30][8]~q ;
wire \Mux23~2_combout ;
wire \Mux23~3_combout ;
wire \Mux23~4_combout ;
wire \Mux23~5_combout ;
wire \Mux23~6_combout ;
wire \Mux23~10_combout ;
wire \Mux23~11_combout ;
wire \Mux23~12_combout ;
wire \Mux23~13_combout ;
wire \Mux23~14_combout ;
wire \Mux23~15_combout ;
wire \Mux23~16_combout ;
wire \Mux23~17_combout ;
wire \Mux23~18_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \Mux24~7_combout ;
wire \Mux24~8_combout ;
wire \Mux24~2_combout ;
wire \Mux24~3_combout ;
wire \Mux24~5_combout ;
wire \Mux24~6_combout ;
wire \rfile[12][7]~q ;
wire \Mux24~17_combout ;
wire \Mux24~18_combout ;
wire \Mux24~10_combout ;
wire \Mux24~11_combout ;
wire \Mux24~14_combout ;
wire \rfile[2][7]~feeder_combout ;
wire \rfile[2][7]~q ;
wire \Mux24~15_combout ;
wire \Mux24~12_combout ;
wire \Mux24~13_combout ;
wire \Mux24~16_combout ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux25~7_combout ;
wire \Mux25~8_combout ;
wire \Mux25~4_combout ;
wire \Mux25~5_combout ;
wire \rfile[26][6]~q ;
wire \Mux25~3_combout ;
wire \Mux25~6_combout ;
wire \rfile[4][6]~q ;
wire \Mux25~10_combout ;
wire \Mux25~11_combout ;
wire \Mux25~14_combout ;
wire \Mux25~15_combout ;
wire \rfile[11][6]~feeder_combout ;
wire \rfile[11][6]~q ;
wire \Mux25~12_combout ;
wire \Mux25~13_combout ;
wire \Mux25~16_combout ;
wire \Mux25~17_combout ;
wire \Mux25~18_combout ;
wire \Mux26~7_combout ;
wire \Mux26~8_combout ;
wire \rfile[22][5]~q ;
wire \rfile[18][5]~feeder_combout ;
wire \rfile[18][5]~q ;
wire \Mux26~2_combout ;
wire \Mux26~3_combout ;
wire \rfile[28][5]~q ;
wire \Mux26~4_combout ;
wire \Mux26~5_combout ;
wire \Mux26~6_combout ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \Mux26~12_combout ;
wire \Mux26~13_combout ;
wire \Mux26~14_combout ;
wire \Mux26~15_combout ;
wire \Mux26~16_combout ;
wire \Mux26~10_combout ;
wire \Mux26~11_combout ;
wire \Mux26~17_combout ;
wire \Mux26~18_combout ;
wire \rfile[19][3]~q ;
wire \Mux60~7_combout ;
wire \Mux60~8_combout ;
wire \Mux60~0_combout ;
wire \Mux60~1_combout ;
wire \Mux60~2_combout ;
wire \Mux60~3_combout ;
wire \rfile[28][3]~q ;
wire \Mux60~4_combout ;
wire \Mux60~5_combout ;
wire \Mux60~6_combout ;
wire \Mux60~12_combout ;
wire \Mux60~13_combout ;
wire \Mux60~14_combout ;
wire \Mux60~15_combout ;
wire \Mux60~16_combout ;
wire \rfile[8][3]~q ;
wire \Mux60~10_combout ;
wire \Mux60~11_combout ;
wire \Mux60~17_combout ;
wire \Mux60~18_combout ;
wire \Mux15~7_combout ;
wire \Mux15~8_combout ;
wire \Mux15~4_combout ;
wire \Mux15~5_combout ;
wire \rfile[22][16]~feeder_combout ;
wire \rfile[22][16]~q ;
wire \rfile[18][16]~q ;
wire \Mux15~2_combout ;
wire \Mux15~3_combout ;
wire \Mux15~6_combout ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \rfile[4][16]~q ;
wire \Mux15~10_combout ;
wire \Mux15~11_combout ;
wire \Mux15~14_combout ;
wire \Mux15~15_combout ;
wire \rfile[8][16]~q ;
wire \Mux15~12_combout ;
wire \Mux15~13_combout ;
wire \Mux15~16_combout ;
wire \Mux15~17_combout ;
wire \Mux15~18_combout ;
wire \Mux16~7_combout ;
wire \Mux16~8_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \rfile[28][15]~feeder_combout ;
wire \rfile[28][15]~q ;
wire \rfile[24][15]~q ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \Mux16~6_combout ;
wire \Mux16~17_combout ;
wire \Mux16~18_combout ;
wire \Mux16~10_combout ;
wire \Mux16~11_combout ;
wire \Mux16~14_combout ;
wire \Mux16~15_combout ;
wire \Mux16~12_combout ;
wire \Mux16~13_combout ;
wire \Mux16~16_combout ;
wire \Mux17~7_combout ;
wire \Mux17~8_combout ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \rfile[24][14]~q ;
wire \Mux17~4_combout ;
wire \Mux17~5_combout ;
wire \Mux17~6_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \Mux17~10_combout ;
wire \Mux17~11_combout ;
wire \Mux17~17_combout ;
wire \Mux17~18_combout ;
wire \Mux17~14_combout ;
wire \Mux17~15_combout ;
wire \Mux17~12_combout ;
wire \Mux17~13_combout ;
wire \Mux17~16_combout ;
wire \Mux18~7_combout ;
wire \Mux18~8_combout ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \rfile[20][13]~feeder_combout ;
wire \rfile[20][13]~q ;
wire \Mux18~4_combout ;
wire \Mux18~5_combout ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \Mux18~6_combout ;
wire \Mux18~17_combout ;
wire \Mux18~18_combout ;
wire \Mux18~14_combout ;
wire \Mux18~15_combout ;
wire \rfile[7][13]~q ;
wire \Mux18~12_combout ;
wire \Mux18~13_combout ;
wire \Mux18~16_combout ;
wire \Mux18~10_combout ;
wire \Mux18~11_combout ;
wire \Mux19~7_combout ;
wire \Mux19~8_combout ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \rfile[30][12]~q ;
wire \Mux19~2_combout ;
wire \Mux19~3_combout ;
wire \Mux19~4_combout ;
wire \rfile[24][12]~q ;
wire \Mux19~5_combout ;
wire \Mux19~6_combout ;
wire \rfile[4][12]~q ;
wire \Mux19~10_combout ;
wire \Mux19~11_combout ;
wire \Mux19~14_combout ;
wire \Mux19~15_combout ;
wire \rfile[10][12]~q ;
wire \rfile[8][12]~q ;
wire \Mux19~12_combout ;
wire \Mux19~13_combout ;
wire \Mux19~16_combout ;
wire \Mux19~17_combout ;
wire \Mux19~18_combout ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \Mux20~7_combout ;
wire \Mux20~8_combout ;
wire \Mux20~4_combout ;
wire \Mux20~5_combout ;
wire \rfile[26][11]~feeder_combout ;
wire \rfile[26][11]~q ;
wire \Mux20~2_combout ;
wire \rfile[30][11]~feeder_combout ;
wire \rfile[30][11]~q ;
wire \Mux20~3_combout ;
wire \Mux20~6_combout ;
wire \Mux20~17_combout ;
wire \Mux20~18_combout ;
wire \Mux20~12_combout ;
wire \rfile[6][11]~feeder_combout ;
wire \rfile[6][11]~q ;
wire \Mux20~13_combout ;
wire \Mux20~14_combout ;
wire \Mux20~15_combout ;
wire \Mux20~16_combout ;
wire \Mux20~10_combout ;
wire \Mux20~11_combout ;
wire \rfile[17][10]~q ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Mux21~7_combout ;
wire \Mux21~8_combout ;
wire \Mux21~5_combout ;
wire \rfile[26][10]~q ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \Mux21~6_combout ;
wire \Mux21~10_combout ;
wire \Mux21~11_combout ;
wire \Mux21~17_combout ;
wire \Mux21~18_combout ;
wire \Mux21~13_combout ;
wire \Mux21~14_combout ;
wire \Mux21~15_combout ;
wire \Mux21~16_combout ;
wire \rfile[20][9]~q ;
wire \Mux22~4_combout ;
wire \Mux22~5_combout ;
wire \Mux22~2_combout ;
wire \Mux22~3_combout ;
wire \Mux22~6_combout ;
wire \Mux22~7_combout ;
wire \Mux22~8_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \Mux22~10_combout ;
wire \Mux22~11_combout ;
wire \rfile[4][9]~q ;
wire \rfile[5][9]~q ;
wire \Mux22~12_combout ;
wire \Mux22~13_combout ;
wire \Mux22~14_combout ;
wire \Mux22~15_combout ;
wire \Mux22~16_combout ;
wire \Mux22~17_combout ;
wire \Mux22~18_combout ;
wire \Mux59~7_combout ;
wire \Mux59~8_combout ;
wire \Mux59~0_combout ;
wire \Mux59~1_combout ;
wire \rfile[30][4]~feeder_combout ;
wire \rfile[30][4]~q ;
wire \Mux59~2_combout ;
wire \Mux59~3_combout ;
wire \Mux59~4_combout ;
wire \Mux59~5_combout ;
wire \Mux59~6_combout ;
wire \Mux59~17_combout ;
wire \Mux59~18_combout ;
wire \Mux59~12_combout ;
wire \Mux59~13_combout ;
wire \Mux59~14_combout ;
wire \Mux59~15_combout ;
wire \Mux59~16_combout ;
wire \Mux59~10_combout ;
wire \Mux59~11_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux0~4_combout ;
wire \rfile[20][31]~q ;
wire \Mux0~5_combout ;
wire \rfile[26][31]~q ;
wire \rfile[18][31]~q ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~6_combout ;
wire \Mux0~7_combout ;
wire \Mux0~8_combout ;
wire \rfile[8][31]~q ;
wire \Mux0~10_combout ;
wire \Mux0~11_combout ;
wire \Mux0~17_combout ;
wire \Mux0~18_combout ;
wire \rfile[7][31]~q ;
wire \rfile[4][31]~q ;
wire \Mux0~12_combout ;
wire \Mux0~13_combout ;
wire \Mux0~15_combout ;
wire \Mux0~16_combout ;
wire \Mux2~7_combout ;
wire \Mux2~8_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \rfile[24][29]~q ;
wire \rfile[16][29]~q ;
wire \Mux2~4_combout ;
wire \Mux2~5_combout ;
wire \Mux2~6_combout ;
wire \Mux2~17_combout ;
wire \Mux2~18_combout ;
wire \Mux2~10_combout ;
wire \Mux2~11_combout ;
wire \rfile[7][29]~q ;
wire \Mux2~12_combout ;
wire \Mux2~13_combout ;
wire \Mux2~14_combout ;
wire \Mux2~15_combout ;
wire \Mux2~16_combout ;
wire \rfile[18][30]~q ;
wire \rfile[22][30]~feeder_combout ;
wire \rfile[22][30]~q ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \Mux1~7_combout ;
wire \Mux1~8_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux1~17_combout ;
wire \Mux1~18_combout ;
wire \rfile[4][30]~q ;
wire \Mux1~10_combout ;
wire \Mux1~11_combout ;
wire \Mux1~14_combout ;
wire \Mux1~15_combout ;
wire \rfile[11][30]~q ;
wire \Mux1~12_combout ;
wire \Mux1~13_combout ;
wire \Mux1~16_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux3~7_combout ;
wire \Mux3~8_combout ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \rfile[28][28]~q ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \Mux3~6_combout ;
wire \Mux3~10_combout ;
wire \Mux3~11_combout ;
wire \Mux3~17_combout ;
wire \Mux3~18_combout ;
wire \Mux3~14_combout ;
wire \Mux3~15_combout ;
wire \Mux3~12_combout ;
wire \Mux3~13_combout ;
wire \Mux3~16_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \rfile[19][27]~q ;
wire \Mux4~7_combout ;
wire \Mux4~8_combout ;
wire \rfile[22][27]~q ;
wire \Mux4~2_combout ;
wire \Mux4~3_combout ;
wire \rfile[28][27]~q ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Mux4~6_combout ;
wire \Mux4~17_combout ;
wire \Mux4~18_combout ;
wire \Mux4~10_combout ;
wire \Mux4~11_combout ;
wire \Mux4~14_combout ;
wire \Mux4~15_combout ;
wire \Mux4~12_combout ;
wire \Mux4~13_combout ;
wire \Mux4~16_combout ;
wire \rfile[17][26]~q ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux5~7_combout ;
wire \Mux5~8_combout ;
wire \rfile[16][26]~q ;
wire \rfile[20][26]~q ;
wire \Mux5~4_combout ;
wire \Mux5~5_combout ;
wire \rfile[18][26]~q ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \Mux5~6_combout ;
wire \Mux5~10_combout ;
wire \Mux5~11_combout ;
wire \Mux5~17_combout ;
wire \Mux5~18_combout ;
wire \Mux5~14_combout ;
wire \Mux5~15_combout ;
wire \rfile[11][26]~q ;
wire \rfile[10][26]~q ;
wire \Mux5~12_combout ;
wire \Mux5~13_combout ;
wire \Mux5~16_combout ;
wire \rfile[19][25]~q ;
wire \Mux6~7_combout ;
wire \Mux6~8_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \rfile[18][25]~q ;
wire \rfile[26][25]~q ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \rfile[28][25]~feeder_combout ;
wire \rfile[28][25]~q ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \Mux6~6_combout ;
wire \Mux6~10_combout ;
wire \Mux6~11_combout ;
wire \Mux6~14_combout ;
wire \Mux6~15_combout ;
wire \Mux6~12_combout ;
wire \Mux6~13_combout ;
wire \Mux6~16_combout ;
wire \Mux6~17_combout ;
wire \Mux6~18_combout ;
wire \Mux7~7_combout ;
wire \Mux7~8_combout ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux7~3_combout ;
wire \rfile[20][24]~q ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \Mux7~6_combout ;
wire \rfile[4][24]~q ;
wire \Mux7~10_combout ;
wire \Mux7~11_combout ;
wire \Mux7~14_combout ;
wire \Mux7~15_combout ;
wire \Mux7~12_combout ;
wire \Mux7~13_combout ;
wire \Mux7~16_combout ;
wire \Mux7~17_combout ;
wire \Mux7~18_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Mux8~7_combout ;
wire \Mux8~8_combout ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \Mux8~6_combout ;
wire \Mux8~17_combout ;
wire \Mux8~18_combout ;
wire \Mux8~14_combout ;
wire \Mux8~15_combout ;
wire \Mux8~12_combout ;
wire \rfile[6][23]~feeder_combout ;
wire \rfile[6][23]~q ;
wire \Mux8~13_combout ;
wire \Mux8~16_combout ;
wire \Mux8~10_combout ;
wire \Mux8~11_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Mux9~7_combout ;
wire \Mux9~8_combout ;
wire \Mux9~2_combout ;
wire \Mux9~3_combout ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux9~6_combout ;
wire \Mux9~17_combout ;
wire \Mux9~18_combout ;
wire \Mux9~10_combout ;
wire \Mux9~11_combout ;
wire \Mux9~14_combout ;
wire \Mux9~15_combout ;
wire \Mux9~12_combout ;
wire \Mux9~13_combout ;
wire \Mux9~16_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \Mux10~7_combout ;
wire \Mux10~8_combout ;
wire \rfile[20][21]~q ;
wire \Mux10~4_combout ;
wire \Mux10~5_combout ;
wire \Mux10~2_combout ;
wire \Mux10~3_combout ;
wire \Mux10~6_combout ;
wire \rfile[4][21]~q ;
wire \Mux10~12_combout ;
wire \Mux10~13_combout ;
wire \Mux10~14_combout ;
wire \Mux10~15_combout ;
wire \Mux10~16_combout ;
wire \Mux10~17_combout ;
wire \Mux10~18_combout ;
wire \Mux10~10_combout ;
wire \Mux10~11_combout ;
wire \Mux11~7_combout ;
wire \Mux11~8_combout ;
wire \rfile[22][20]~q ;
wire \Mux11~2_combout ;
wire \Mux11~3_combout ;
wire \rfile[24][20]~q ;
wire \Mux11~4_combout ;
wire \Mux11~5_combout ;
wire \Mux11~6_combout ;
wire \rfile[25][20]~q ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \rfile[1][20]~q ;
wire \Mux11~14_combout ;
wire \Mux11~15_combout ;
wire \Mux11~12_combout ;
wire \rfile[11][20]~q ;
wire \Mux11~13_combout ;
wire \Mux11~16_combout ;
wire \Mux11~17_combout ;
wire \Mux11~18_combout ;
wire \Mux11~10_combout ;
wire \Mux11~11_combout ;
wire \Mux12~7_combout ;
wire \Mux12~8_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \Mux12~4_combout ;
wire \Mux12~5_combout ;
wire \Mux12~6_combout ;
wire \Mux12~17_combout ;
wire \Mux12~18_combout ;
wire \Mux12~10_combout ;
wire \Mux12~11_combout ;
wire \rfile[4][19]~q ;
wire \rfile[5][19]~q ;
wire \Mux12~12_combout ;
wire \Mux12~13_combout ;
wire \Mux12~14_combout ;
wire \Mux12~15_combout ;
wire \Mux12~16_combout ;
wire \Mux13~7_combout ;
wire \Mux13~8_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \Mux13~4_combout ;
wire \Mux13~5_combout ;
wire \Mux13~6_combout ;
wire \Mux13~10_combout ;
wire \Mux13~11_combout ;
wire \Mux13~17_combout ;
wire \Mux13~18_combout ;
wire \Mux13~14_combout ;
wire \Mux13~15_combout ;
wire \Mux13~12_combout ;
wire \Mux13~13_combout ;
wire \Mux13~16_combout ;
wire \rfile[20][17]~feeder_combout ;
wire \rfile[20][17]~q ;
wire \Mux14~4_combout ;
wire \Mux14~5_combout ;
wire \rfile[22][17]~q ;
wire \Mux14~3_combout ;
wire \Mux14~6_combout ;
wire \Mux14~7_combout ;
wire \Mux14~8_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \Mux14~10_combout ;
wire \Mux14~11_combout ;
wire \Mux14~12_combout ;
wire \Mux14~13_combout ;
wire \Mux14~14_combout ;
wire \Mux14~15_combout ;
wire \Mux14~16_combout ;
wire \Mux14~17_combout ;
wire \Mux14~18_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux31~7_combout ;
wire \Mux31~8_combout ;
wire \Mux31~4_combout ;
wire \rfile[28][0]~q ;
wire \Mux31~5_combout ;
wire \Mux31~2_combout ;
wire \Mux31~3_combout ;
wire \Mux31~6_combout ;
wire \Mux31~10_combout ;
wire \Mux31~11_combout ;
wire \rfile[12][0]~q ;
wire \Mux31~17_combout ;
wire \Mux31~18_combout ;
wire \Mux31~14_combout ;
wire \Mux31~15_combout ;
wire \Mux31~12_combout ;
wire \Mux31~13_combout ;
wire \Mux31~16_combout ;


// Location: LCCOMB_X75_Y34_N22
cycloneive_lcell_comb \Mux32~2 (
// Equation(s):
// \Mux32~2_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[26][31]~q )) # (!instruction_D[19] & ((\rfile[18][31]~q )))))

	.dataa(\rfile[26][31]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[18][31]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~2 .lut_mask = 16'hEE30;
defparam \Mux32~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N12
cycloneive_lcell_comb \Mux33~2 (
// Equation(s):
// \Mux33~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[22][30]~q ))) # (!instruction_D[18] & (\rfile[18][30]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][30]~q ),
	.datad(\rfile[22][30]~q ),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~2 .lut_mask = 16'hDC98;
defparam \Mux33~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N27
dffeas \rfile[28][30] (
	.clk(!CLK),
	.d(\rfile[28][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][30] .is_wysiwyg = "true";
defparam \rfile[28][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N22
cycloneive_lcell_comb \Mux34~4 (
// Equation(s):
// \Mux34~4_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[24][29]~q ))) # (!instruction_D[19] & (\rfile[16][29]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[16][29]~q ),
	.datad(\rfile[24][29]~q ),
	.cin(gnd),
	.combout(\Mux34~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~4 .lut_mask = 16'hDC98;
defparam \Mux34~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N31
dffeas \rfile[7][27] (
	.clk(!CLK),
	.d(\rfile[7][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][27] .is_wysiwyg = "true";
defparam \rfile[7][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N20
cycloneive_lcell_comb \Mux37~4 (
// Equation(s):
// \Mux37~4_combout  = (instruction_D[19] & (((instruction_D[18])))) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[20][26]~q ))) # (!instruction_D[18] & (\rfile[16][26]~q ))))

	.dataa(\rfile[16][26]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[20][26]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux37~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~4 .lut_mask = 16'hFC22;
defparam \Mux37~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N0
cycloneive_lcell_comb \Mux38~2 (
// Equation(s):
// \Mux38~2_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[26][25]~q )) # (!instruction_D[19] & ((\rfile[18][25]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[26][25]~q ),
	.datad(\rfile[18][25]~q ),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~2 .lut_mask = 16'hD9C8;
defparam \Mux38~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y31_N31
dffeas \rfile[16][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][24] .is_wysiwyg = "true";
defparam \rfile[16][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N30
cycloneive_lcell_comb \Mux39~4 (
// Equation(s):
// \Mux39~4_combout  = (instruction_D[19] & (((instruction_D[18])))) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[20][24]~q )) # (!instruction_D[18] & ((\rfile[16][24]~q )))))

	.dataa(instruction_D_19),
	.datab(\rfile[20][24]~q ),
	.datac(\rfile[16][24]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux39~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~4 .lut_mask = 16'hEE50;
defparam \Mux39~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N1
dffeas \rfile[9][24] (
	.clk(!CLK),
	.d(\rfile[9][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][24] .is_wysiwyg = "true";
defparam \rfile[9][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y30_N11
dffeas \rfile[28][22] (
	.clk(!CLK),
	.d(\rfile[28][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][22] .is_wysiwyg = "true";
defparam \rfile[28][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N2
cycloneive_lcell_comb \Mux44~12 (
// Equation(s):
// \Mux44~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[5][19]~q )) # (!instruction_D[16] & ((\rfile[4][19]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[5][19]~q ),
	.datad(\rfile[4][19]~q ),
	.cin(gnd),
	.combout(\Mux44~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~12 .lut_mask = 16'hD9C8;
defparam \Mux44~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N31
dffeas \rfile[5][18] (
	.clk(!CLK),
	.d(\rfile[5][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][18] .is_wysiwyg = "true";
defparam \rfile[5][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N30
cycloneive_lcell_comb \Mux47~2 (
// Equation(s):
// \Mux47~2_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[22][16]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[18][16]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[18][16]~q ),
	.datad(\rfile[22][16]~q ),
	.cin(gnd),
	.combout(\Mux47~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~2 .lut_mask = 16'hBA98;
defparam \Mux47~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y30_N31
dffeas \rfile[24][16] (
	.clk(!CLK),
	.d(\rfile[24][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][16] .is_wysiwyg = "true";
defparam \rfile[24][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N4
cycloneive_lcell_comb \Mux51~12 (
// Equation(s):
// \Mux51~12_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][12]~q ))) # (!instruction_D[17] & (\rfile[8][12]~q ))))

	.dataa(instruction_D_16),
	.datab(\rfile[8][12]~q ),
	.datac(\rfile[10][12]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux51~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~12 .lut_mask = 16'hFA44;
defparam \Mux51~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N26
cycloneive_lcell_comb \Mux54~12 (
// Equation(s):
// \Mux54~12_combout  = (instruction_D[16] & (((\rfile[5][9]~q ) # (instruction_D[17])))) # (!instruction_D[16] & (\rfile[4][9]~q  & ((!instruction_D[17]))))

	.dataa(\rfile[4][9]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[5][9]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux54~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~12 .lut_mask = 16'hCCE2;
defparam \Mux54~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y27_N13
dffeas \rfile[2][9] (
	.clk(!CLK),
	.d(\rfile[2][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][9] .is_wysiwyg = "true";
defparam \rfile[2][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y30_N13
dffeas \rfile[28][8] (
	.clk(!CLK),
	.d(\rfile[28][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][8] .is_wysiwyg = "true";
defparam \rfile[28][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y29_N31
dffeas \rfile[6][7] (
	.clk(!CLK),
	.d(\rfile[6][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][7] .is_wysiwyg = "true";
defparam \rfile[6][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N17
dffeas \rfile[26][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][1] .is_wysiwyg = "true";
defparam \rfile[26][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N11
dffeas \rfile[18][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][1] .is_wysiwyg = "true";
defparam \rfile[18][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N10
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\rfile[26][1]~q ))) # (!instruction_D[24] & (\rfile[18][1]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[18][1]~q ),
	.datad(\rfile[26][1]~q ),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'hDC98;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N31
dffeas \rfile[4][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][1] .is_wysiwyg = "true";
defparam \rfile[4][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N30
cycloneive_lcell_comb \Mux30~12 (
// Equation(s):
// \Mux30~12_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[5][1]~q )) # (!instruction_D[21] & ((\rfile[4][1]~q )))))

	.dataa(instruction_D_22),
	.datab(\rfile[5][1]~q ),
	.datac(\rfile[4][1]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux30~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~12 .lut_mask = 16'hEE50;
defparam \Mux30~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N11
dffeas \rfile[2][1] (
	.clk(!CLK),
	.d(\rfile[2][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][1] .is_wysiwyg = "true";
defparam \rfile[2][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N7
dffeas \rfile[12][1] (
	.clk(!CLK),
	.d(\rfile[12][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][1] .is_wysiwyg = "true";
defparam \rfile[12][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N16
cycloneive_lcell_comb \Mux62~2 (
// Equation(s):
// \Mux62~2_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[26][1]~q )) # (!instruction_D[19] & ((\rfile[18][1]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[26][1]~q ),
	.datad(\rfile[18][1]~q ),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~2 .lut_mask = 16'hD9C8;
defparam \Mux62~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N10
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[24][7]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[16][7]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[24][7]~q ),
	.datad(\rfile[16][7]~q ),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'hB9A8;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N26
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[22][6]~q )))) # (!instruction_D[23] & (!instruction_D[24] & (\rfile[18][6]~q )))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[18][6]~q ),
	.datad(\rfile[22][6]~q ),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'hBA98;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N26
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[20][10]~q ))) # (!instruction_D[23] & (\rfile[16][10]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[16][10]~q ),
	.datad(\rfile[20][10]~q ),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hDC98;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N28
cycloneive_lcell_comb \Mux21~12 (
// Equation(s):
// \Mux21~12_combout  = (instruction_D[22] & (((\rfile[10][10]~q ) # (instruction_D[21])))) # (!instruction_D[22] & (\rfile[8][10]~q  & ((!instruction_D[21]))))

	.dataa(\rfile[8][10]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[10][10]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux21~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~12 .lut_mask = 16'hCCE2;
defparam \Mux21~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N14
cycloneive_lcell_comb \Mux0~14 (
// Equation(s):
// \Mux0~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][31]~q ))) # (!instruction_D[22] & (\rfile[1][31]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][31]~q ),
	.datad(\rfile[3][31]~q ),
	.cin(gnd),
	.combout(\Mux0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~14 .lut_mask = 16'hC840;
defparam \Mux0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N30
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[22][24]~q )) # (!instruction_D[23] & ((\rfile[18][24]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[22][24]~q ),
	.datad(\rfile[18][24]~q ),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hD9C8;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N14
cycloneive_lcell_comb \Mux14~2 (
// Equation(s):
// \Mux14~2_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\rfile[26][17]~q ))) # (!instruction_D[24] & (\rfile[18][17]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[18][17]~q ),
	.datad(\rfile[26][17]~q ),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~2 .lut_mask = 16'hDC98;
defparam \Mux14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N26
cycloneive_lcell_comb \rfile[28][30]~feeder (
// Equation(s):
// \rfile[28][30]~feeder_combout  = \wdat_WB[30]~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_30),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[28][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][30]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[28][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N30
cycloneive_lcell_comb \rfile[7][27]~feeder (
// Equation(s):
// \rfile[7][27]~feeder_combout  = \wdat_WB[27]~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_27),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[7][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[7][27]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[7][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N0
cycloneive_lcell_comb \rfile[9][24]~feeder (
// Equation(s):
// \rfile[9][24]~feeder_combout  = \wdat_WB[24]~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_24),
	.cin(gnd),
	.combout(\rfile[9][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][24]~feeder .lut_mask = 16'hFF00;
defparam \rfile[9][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N10
cycloneive_lcell_comb \rfile[28][22]~feeder (
// Equation(s):
// \rfile[28][22]~feeder_combout  = \wdat_WB[22]~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[28][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][22]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[28][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N30
cycloneive_lcell_comb \rfile[5][18]~feeder (
// Equation(s):
// \rfile[5][18]~feeder_combout  = \wdat_WB[18]~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_18),
	.cin(gnd),
	.combout(\rfile[5][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[5][18]~feeder .lut_mask = 16'hFF00;
defparam \rfile[5][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N30
cycloneive_lcell_comb \rfile[24][16]~feeder (
// Equation(s):
// \rfile[24][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_16),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[24][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[24][16]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[24][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N12
cycloneive_lcell_comb \rfile[2][9]~feeder (
// Equation(s):
// \rfile[2][9]~feeder_combout  = \wdat_WB[9]~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_9),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[2][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][9]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[2][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N12
cycloneive_lcell_comb \rfile[28][8]~feeder (
// Equation(s):
// \rfile[28][8]~feeder_combout  = \wdat_WB[8]~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[28][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][8]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[28][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N30
cycloneive_lcell_comb \rfile[6][7]~feeder (
// Equation(s):
// \rfile[6][7]~feeder_combout  = \wdat_WB[7]~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[6][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][7]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[6][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N10
cycloneive_lcell_comb \rfile[2][1]~feeder (
// Equation(s):
// \rfile[2][1]~feeder_combout  = \wdat_WB[1]~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_1),
	.cin(gnd),
	.combout(\rfile[2][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][1]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N6
cycloneive_lcell_comb \rfile[12][1]~feeder (
// Equation(s):
// \rfile[12][1]~feeder_combout  = \wdat_WB[1]~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_1),
	.cin(gnd),
	.combout(\rfile[12][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[12][1]~feeder .lut_mask = 16'hFF00;
defparam \rfile[12][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N16
cycloneive_lcell_comb \Mux32~9 (
// Equation(s):
// Mux32 = (instruction_D[16] & ((\Mux32~6_combout  & ((\Mux32~8_combout ))) # (!\Mux32~6_combout  & (\Mux32~1_combout )))) # (!instruction_D[16] & (((\Mux32~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux32~1_combout ),
	.datac(\Mux32~8_combout ),
	.datad(\Mux32~6_combout ),
	.cin(gnd),
	.combout(Mux32),
	.cout());
// synopsys translate_off
defparam \Mux32~9 .lut_mask = 16'hF588;
defparam \Mux32~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N18
cycloneive_lcell_comb \Mux32~19 (
// Equation(s):
// Mux321 = (instruction_D[19] & ((\Mux32~16_combout  & ((\Mux32~18_combout ))) # (!\Mux32~16_combout  & (\Mux32~11_combout )))) # (!instruction_D[19] & (((\Mux32~16_combout ))))

	.dataa(instruction_D_19),
	.datab(\Mux32~11_combout ),
	.datac(\Mux32~16_combout ),
	.datad(\Mux32~18_combout ),
	.cin(gnd),
	.combout(Mux321),
	.cout());
// synopsys translate_off
defparam \Mux32~19 .lut_mask = 16'hF858;
defparam \Mux32~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N10
cycloneive_lcell_comb \Mux33~9 (
// Equation(s):
// Mux33 = (instruction_D[16] & ((\Mux33~6_combout  & ((\Mux33~8_combout ))) # (!\Mux33~6_combout  & (\Mux33~1_combout )))) # (!instruction_D[16] & (((\Mux33~6_combout ))))

	.dataa(\Mux33~1_combout ),
	.datab(instruction_D_16),
	.datac(\Mux33~8_combout ),
	.datad(\Mux33~6_combout ),
	.cin(gnd),
	.combout(Mux33),
	.cout());
// synopsys translate_off
defparam \Mux33~9 .lut_mask = 16'hF388;
defparam \Mux33~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N16
cycloneive_lcell_comb \Mux33~19 (
// Equation(s):
// Mux331 = (instruction_D[18] & ((\Mux33~16_combout  & (\Mux33~18_combout )) # (!\Mux33~16_combout  & ((\Mux33~11_combout ))))) # (!instruction_D[18] & (((\Mux33~16_combout ))))

	.dataa(\Mux33~18_combout ),
	.datab(instruction_D_18),
	.datac(\Mux33~16_combout ),
	.datad(\Mux33~11_combout ),
	.cin(gnd),
	.combout(Mux331),
	.cout());
// synopsys translate_off
defparam \Mux33~19 .lut_mask = 16'hBCB0;
defparam \Mux33~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N30
cycloneive_lcell_comb \Mux34~9 (
// Equation(s):
// Mux34 = (instruction_D[16] & ((\Mux34~6_combout  & ((\Mux34~8_combout ))) # (!\Mux34~6_combout  & (\Mux34~1_combout )))) # (!instruction_D[16] & (((\Mux34~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux34~1_combout ),
	.datac(\Mux34~6_combout ),
	.datad(\Mux34~8_combout ),
	.cin(gnd),
	.combout(Mux34),
	.cout());
// synopsys translate_off
defparam \Mux34~9 .lut_mask = 16'hF858;
defparam \Mux34~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N24
cycloneive_lcell_comb \Mux34~19 (
// Equation(s):
// Mux341 = (instruction_D[19] & ((\Mux34~16_combout  & ((\Mux34~18_combout ))) # (!\Mux34~16_combout  & (\Mux34~11_combout )))) # (!instruction_D[19] & (((\Mux34~16_combout ))))

	.dataa(instruction_D_19),
	.datab(\Mux34~11_combout ),
	.datac(\Mux34~18_combout ),
	.datad(\Mux34~16_combout ),
	.cin(gnd),
	.combout(Mux341),
	.cout());
// synopsys translate_off
defparam \Mux34~19 .lut_mask = 16'hF588;
defparam \Mux34~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N30
cycloneive_lcell_comb \Mux35~9 (
// Equation(s):
// Mux35 = (instruction_D[16] & ((\Mux35~6_combout  & (\Mux35~8_combout )) # (!\Mux35~6_combout  & ((\Mux35~1_combout ))))) # (!instruction_D[16] & (((\Mux35~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux35~8_combout ),
	.datac(\Mux35~6_combout ),
	.datad(\Mux35~1_combout ),
	.cin(gnd),
	.combout(Mux35),
	.cout());
// synopsys translate_off
defparam \Mux35~9 .lut_mask = 16'hDAD0;
defparam \Mux35~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N4
cycloneive_lcell_comb \Mux35~19 (
// Equation(s):
// Mux351 = (instruction_D[18] & ((\Mux35~16_combout  & (\Mux35~18_combout )) # (!\Mux35~16_combout  & ((\Mux35~11_combout ))))) # (!instruction_D[18] & (((\Mux35~16_combout ))))

	.dataa(\Mux35~18_combout ),
	.datab(instruction_D_18),
	.datac(\Mux35~16_combout ),
	.datad(\Mux35~11_combout ),
	.cin(gnd),
	.combout(Mux351),
	.cout());
// synopsys translate_off
defparam \Mux35~19 .lut_mask = 16'hBCB0;
defparam \Mux35~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N8
cycloneive_lcell_comb \Mux36~9 (
// Equation(s):
// Mux36 = (instruction_D[16] & ((\Mux36~6_combout  & (\Mux36~8_combout )) # (!\Mux36~6_combout  & ((\Mux36~1_combout ))))) # (!instruction_D[16] & (((\Mux36~6_combout ))))

	.dataa(\Mux36~8_combout ),
	.datab(instruction_D_16),
	.datac(\Mux36~1_combout ),
	.datad(\Mux36~6_combout ),
	.cin(gnd),
	.combout(Mux36),
	.cout());
// synopsys translate_off
defparam \Mux36~9 .lut_mask = 16'hBBC0;
defparam \Mux36~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N16
cycloneive_lcell_comb \Mux36~19 (
// Equation(s):
// Mux361 = (instruction_D[19] & ((\Mux36~16_combout  & (\Mux36~18_combout )) # (!\Mux36~16_combout  & ((\Mux36~11_combout ))))) # (!instruction_D[19] & (((\Mux36~16_combout ))))

	.dataa(instruction_D_19),
	.datab(\Mux36~18_combout ),
	.datac(\Mux36~16_combout ),
	.datad(\Mux36~11_combout ),
	.cin(gnd),
	.combout(Mux361),
	.cout());
// synopsys translate_off
defparam \Mux36~19 .lut_mask = 16'hDAD0;
defparam \Mux36~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N16
cycloneive_lcell_comb \Mux37~9 (
// Equation(s):
// Mux37 = (instruction_D[16] & ((\Mux37~6_combout  & (\Mux37~8_combout )) # (!\Mux37~6_combout  & ((\Mux37~1_combout ))))) # (!instruction_D[16] & (((\Mux37~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux37~8_combout ),
	.datac(\Mux37~6_combout ),
	.datad(\Mux37~1_combout ),
	.cin(gnd),
	.combout(Mux37),
	.cout());
// synopsys translate_off
defparam \Mux37~9 .lut_mask = 16'hDAD0;
defparam \Mux37~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N4
cycloneive_lcell_comb \Mux37~19 (
// Equation(s):
// Mux371 = (\Mux37~16_combout  & (((\Mux37~18_combout )) # (!instruction_D[18]))) # (!\Mux37~16_combout  & (instruction_D[18] & (\Mux37~11_combout )))

	.dataa(\Mux37~16_combout ),
	.datab(instruction_D_18),
	.datac(\Mux37~11_combout ),
	.datad(\Mux37~18_combout ),
	.cin(gnd),
	.combout(Mux371),
	.cout());
// synopsys translate_off
defparam \Mux37~19 .lut_mask = 16'hEA62;
defparam \Mux37~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N22
cycloneive_lcell_comb \Mux38~9 (
// Equation(s):
// Mux38 = (instruction_D[16] & ((\Mux38~6_combout  & (\Mux38~8_combout )) # (!\Mux38~6_combout  & ((\Mux38~1_combout ))))) # (!instruction_D[16] & (((\Mux38~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux38~8_combout ),
	.datac(\Mux38~1_combout ),
	.datad(\Mux38~6_combout ),
	.cin(gnd),
	.combout(Mux38),
	.cout());
// synopsys translate_off
defparam \Mux38~9 .lut_mask = 16'hDDA0;
defparam \Mux38~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N26
cycloneive_lcell_comb \Mux38~19 (
// Equation(s):
// Mux381 = (instruction_D[19] & ((\Mux38~16_combout  & (\Mux38~18_combout )) # (!\Mux38~16_combout  & ((\Mux38~11_combout ))))) # (!instruction_D[19] & (((\Mux38~16_combout ))))

	.dataa(\Mux38~18_combout ),
	.datab(instruction_D_19),
	.datac(\Mux38~11_combout ),
	.datad(\Mux38~16_combout ),
	.cin(gnd),
	.combout(Mux381),
	.cout());
// synopsys translate_off
defparam \Mux38~19 .lut_mask = 16'hBBC0;
defparam \Mux38~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N14
cycloneive_lcell_comb \Mux39~9 (
// Equation(s):
// Mux39 = (instruction_D[16] & ((\Mux39~6_combout  & ((\Mux39~8_combout ))) # (!\Mux39~6_combout  & (\Mux39~1_combout )))) # (!instruction_D[16] & (((\Mux39~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux39~1_combout ),
	.datac(\Mux39~6_combout ),
	.datad(\Mux39~8_combout ),
	.cin(gnd),
	.combout(Mux39),
	.cout());
// synopsys translate_off
defparam \Mux39~9 .lut_mask = 16'hF858;
defparam \Mux39~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N24
cycloneive_lcell_comb \Mux39~19 (
// Equation(s):
// Mux391 = (instruction_D[18] & ((\Mux39~16_combout  & ((\Mux39~18_combout ))) # (!\Mux39~16_combout  & (\Mux39~11_combout )))) # (!instruction_D[18] & (((\Mux39~16_combout ))))

	.dataa(instruction_D_18),
	.datab(\Mux39~11_combout ),
	.datac(\Mux39~16_combout ),
	.datad(\Mux39~18_combout ),
	.cin(gnd),
	.combout(Mux391),
	.cout());
// synopsys translate_off
defparam \Mux39~19 .lut_mask = 16'hF858;
defparam \Mux39~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N2
cycloneive_lcell_comb \Mux40~9 (
// Equation(s):
// Mux40 = (instruction_D[16] & ((\Mux40~6_combout  & ((\Mux40~8_combout ))) # (!\Mux40~6_combout  & (\Mux40~1_combout )))) # (!instruction_D[16] & (((\Mux40~6_combout ))))

	.dataa(\Mux40~1_combout ),
	.datab(instruction_D_16),
	.datac(\Mux40~8_combout ),
	.datad(\Mux40~6_combout ),
	.cin(gnd),
	.combout(Mux40),
	.cout());
// synopsys translate_off
defparam \Mux40~9 .lut_mask = 16'hF388;
defparam \Mux40~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N18
cycloneive_lcell_comb \Mux40~19 (
// Equation(s):
// Mux401 = (instruction_D[19] & ((\Mux40~16_combout  & ((\Mux40~18_combout ))) # (!\Mux40~16_combout  & (\Mux40~11_combout )))) # (!instruction_D[19] & (\Mux40~16_combout ))

	.dataa(instruction_D_19),
	.datab(\Mux40~16_combout ),
	.datac(\Mux40~11_combout ),
	.datad(\Mux40~18_combout ),
	.cin(gnd),
	.combout(Mux401),
	.cout());
// synopsys translate_off
defparam \Mux40~19 .lut_mask = 16'hEC64;
defparam \Mux40~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N6
cycloneive_lcell_comb \Mux41~9 (
// Equation(s):
// Mux41 = (instruction_D[16] & ((\Mux41~6_combout  & ((\Mux41~8_combout ))) # (!\Mux41~6_combout  & (\Mux41~1_combout )))) # (!instruction_D[16] & (((\Mux41~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux41~1_combout ),
	.datac(\Mux41~8_combout ),
	.datad(\Mux41~6_combout ),
	.cin(gnd),
	.combout(Mux41),
	.cout());
// synopsys translate_off
defparam \Mux41~9 .lut_mask = 16'hF588;
defparam \Mux41~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N26
cycloneive_lcell_comb \Mux41~19 (
// Equation(s):
// Mux411 = (instruction_D[18] & ((\Mux41~16_combout  & (\Mux41~18_combout )) # (!\Mux41~16_combout  & ((\Mux41~11_combout ))))) # (!instruction_D[18] & (((\Mux41~16_combout ))))

	.dataa(\Mux41~18_combout ),
	.datab(instruction_D_18),
	.datac(\Mux41~16_combout ),
	.datad(\Mux41~11_combout ),
	.cin(gnd),
	.combout(Mux411),
	.cout());
// synopsys translate_off
defparam \Mux41~19 .lut_mask = 16'hBCB0;
defparam \Mux41~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N6
cycloneive_lcell_comb \Mux42~9 (
// Equation(s):
// Mux42 = (instruction_D[16] & ((\Mux42~6_combout  & ((\Mux42~8_combout ))) # (!\Mux42~6_combout  & (\Mux42~1_combout )))) # (!instruction_D[16] & (((\Mux42~6_combout ))))

	.dataa(\Mux42~1_combout ),
	.datab(instruction_D_16),
	.datac(\Mux42~8_combout ),
	.datad(\Mux42~6_combout ),
	.cin(gnd),
	.combout(Mux42),
	.cout());
// synopsys translate_off
defparam \Mux42~9 .lut_mask = 16'hF388;
defparam \Mux42~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N18
cycloneive_lcell_comb \Mux42~19 (
// Equation(s):
// Mux421 = (instruction_D[19] & ((\Mux42~16_combout  & (\Mux42~18_combout )) # (!\Mux42~16_combout  & ((\Mux42~11_combout ))))) # (!instruction_D[19] & (((\Mux42~16_combout ))))

	.dataa(\Mux42~18_combout ),
	.datab(instruction_D_19),
	.datac(\Mux42~11_combout ),
	.datad(\Mux42~16_combout ),
	.cin(gnd),
	.combout(Mux421),
	.cout());
// synopsys translate_off
defparam \Mux42~19 .lut_mask = 16'hBBC0;
defparam \Mux42~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N4
cycloneive_lcell_comb \Mux43~9 (
// Equation(s):
// Mux43 = (instruction_D[16] & ((\Mux43~6_combout  & ((\Mux43~8_combout ))) # (!\Mux43~6_combout  & (\Mux43~1_combout )))) # (!instruction_D[16] & (((\Mux43~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux43~1_combout ),
	.datac(\Mux43~6_combout ),
	.datad(\Mux43~8_combout ),
	.cin(gnd),
	.combout(Mux43),
	.cout());
// synopsys translate_off
defparam \Mux43~9 .lut_mask = 16'hF858;
defparam \Mux43~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N10
cycloneive_lcell_comb \Mux43~19 (
// Equation(s):
// Mux431 = (\Mux43~16_combout  & ((\Mux43~18_combout ) # ((!instruction_D[18])))) # (!\Mux43~16_combout  & (((instruction_D[18] & \Mux43~11_combout ))))

	.dataa(\Mux43~18_combout ),
	.datab(\Mux43~16_combout ),
	.datac(instruction_D_18),
	.datad(\Mux43~11_combout ),
	.cin(gnd),
	.combout(Mux431),
	.cout());
// synopsys translate_off
defparam \Mux43~19 .lut_mask = 16'hBC8C;
defparam \Mux43~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N8
cycloneive_lcell_comb \Mux44~9 (
// Equation(s):
// Mux44 = (instruction_D[16] & ((\Mux44~6_combout  & ((\Mux44~8_combout ))) # (!\Mux44~6_combout  & (\Mux44~1_combout )))) # (!instruction_D[16] & (((\Mux44~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux44~1_combout ),
	.datac(\Mux44~8_combout ),
	.datad(\Mux44~6_combout ),
	.cin(gnd),
	.combout(Mux44),
	.cout());
// synopsys translate_off
defparam \Mux44~9 .lut_mask = 16'hF588;
defparam \Mux44~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N12
cycloneive_lcell_comb \Mux44~19 (
// Equation(s):
// Mux441 = (instruction_D[19] & ((\Mux44~16_combout  & ((\Mux44~18_combout ))) # (!\Mux44~16_combout  & (\Mux44~11_combout )))) # (!instruction_D[19] & (((\Mux44~16_combout ))))

	.dataa(instruction_D_19),
	.datab(\Mux44~11_combout ),
	.datac(\Mux44~16_combout ),
	.datad(\Mux44~18_combout ),
	.cin(gnd),
	.combout(Mux441),
	.cout());
// synopsys translate_off
defparam \Mux44~19 .lut_mask = 16'hF858;
defparam \Mux44~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N26
cycloneive_lcell_comb \Mux45~9 (
// Equation(s):
// Mux45 = (instruction_D[16] & ((\Mux45~6_combout  & ((\Mux45~8_combout ))) # (!\Mux45~6_combout  & (\Mux45~1_combout )))) # (!instruction_D[16] & (((\Mux45~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux45~1_combout ),
	.datac(\Mux45~8_combout ),
	.datad(\Mux45~6_combout ),
	.cin(gnd),
	.combout(Mux45),
	.cout());
// synopsys translate_off
defparam \Mux45~9 .lut_mask = 16'hF588;
defparam \Mux45~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N12
cycloneive_lcell_comb \Mux45~19 (
// Equation(s):
// Mux451 = (instruction_D[18] & ((\Mux45~16_combout  & ((\Mux45~18_combout ))) # (!\Mux45~16_combout  & (\Mux45~11_combout )))) # (!instruction_D[18] & (((\Mux45~16_combout ))))

	.dataa(\Mux45~11_combout ),
	.datab(instruction_D_18),
	.datac(\Mux45~18_combout ),
	.datad(\Mux45~16_combout ),
	.cin(gnd),
	.combout(Mux451),
	.cout());
// synopsys translate_off
defparam \Mux45~19 .lut_mask = 16'hF388;
defparam \Mux45~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N6
cycloneive_lcell_comb \Mux46~9 (
// Equation(s):
// Mux46 = (\Mux46~6_combout  & (((\Mux46~8_combout )) # (!instruction_D[16]))) # (!\Mux46~6_combout  & (instruction_D[16] & ((\Mux46~1_combout ))))

	.dataa(\Mux46~6_combout ),
	.datab(instruction_D_16),
	.datac(\Mux46~8_combout ),
	.datad(\Mux46~1_combout ),
	.cin(gnd),
	.combout(Mux46),
	.cout());
// synopsys translate_off
defparam \Mux46~9 .lut_mask = 16'hE6A2;
defparam \Mux46~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N30
cycloneive_lcell_comb \Mux46~19 (
// Equation(s):
// Mux461 = (instruction_D[19] & ((\Mux46~16_combout  & ((\Mux46~18_combout ))) # (!\Mux46~16_combout  & (\Mux46~11_combout )))) # (!instruction_D[19] & (\Mux46~16_combout ))

	.dataa(instruction_D_19),
	.datab(\Mux46~16_combout ),
	.datac(\Mux46~11_combout ),
	.datad(\Mux46~18_combout ),
	.cin(gnd),
	.combout(Mux461),
	.cout());
// synopsys translate_off
defparam \Mux46~19 .lut_mask = 16'hEC64;
defparam \Mux46~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N6
cycloneive_lcell_comb \Mux47~9 (
// Equation(s):
// Mux47 = (instruction_D[16] & ((\Mux47~6_combout  & (\Mux47~8_combout )) # (!\Mux47~6_combout  & ((\Mux47~1_combout ))))) # (!instruction_D[16] & (((\Mux47~6_combout ))))

	.dataa(\Mux47~8_combout ),
	.datab(instruction_D_16),
	.datac(\Mux47~6_combout ),
	.datad(\Mux47~1_combout ),
	.cin(gnd),
	.combout(Mux47),
	.cout());
// synopsys translate_off
defparam \Mux47~9 .lut_mask = 16'hBCB0;
defparam \Mux47~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N0
cycloneive_lcell_comb \Mux47~19 (
// Equation(s):
// Mux471 = (\Mux47~16_combout  & (((\Mux47~18_combout )) # (!instruction_D[18]))) # (!\Mux47~16_combout  & (instruction_D[18] & (\Mux47~11_combout )))

	.dataa(\Mux47~16_combout ),
	.datab(instruction_D_18),
	.datac(\Mux47~11_combout ),
	.datad(\Mux47~18_combout ),
	.cin(gnd),
	.combout(Mux471),
	.cout());
// synopsys translate_off
defparam \Mux47~19 .lut_mask = 16'hEA62;
defparam \Mux47~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N14
cycloneive_lcell_comb \Mux48~9 (
// Equation(s):
// Mux48 = (instruction_D[16] & ((\Mux48~6_combout  & ((\Mux48~8_combout ))) # (!\Mux48~6_combout  & (\Mux48~1_combout )))) # (!instruction_D[16] & (((\Mux48~6_combout ))))

	.dataa(\Mux48~1_combout ),
	.datab(instruction_D_16),
	.datac(\Mux48~8_combout ),
	.datad(\Mux48~6_combout ),
	.cin(gnd),
	.combout(Mux48),
	.cout());
// synopsys translate_off
defparam \Mux48~9 .lut_mask = 16'hF388;
defparam \Mux48~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N18
cycloneive_lcell_comb \Mux48~19 (
// Equation(s):
// Mux481 = (instruction_D[19] & ((\Mux48~16_combout  & (\Mux48~18_combout )) # (!\Mux48~16_combout  & ((\Mux48~11_combout ))))) # (!instruction_D[19] & (((\Mux48~16_combout ))))

	.dataa(\Mux48~18_combout ),
	.datab(instruction_D_19),
	.datac(\Mux48~11_combout ),
	.datad(\Mux48~16_combout ),
	.cin(gnd),
	.combout(Mux481),
	.cout());
// synopsys translate_off
defparam \Mux48~19 .lut_mask = 16'hBBC0;
defparam \Mux48~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N4
cycloneive_lcell_comb \Mux49~9 (
// Equation(s):
// Mux49 = (instruction_D[16] & ((\Mux49~6_combout  & (\Mux49~8_combout )) # (!\Mux49~6_combout  & ((\Mux49~1_combout ))))) # (!instruction_D[16] & (((\Mux49~6_combout ))))

	.dataa(\Mux49~8_combout ),
	.datab(instruction_D_16),
	.datac(\Mux49~6_combout ),
	.datad(\Mux49~1_combout ),
	.cin(gnd),
	.combout(Mux49),
	.cout());
// synopsys translate_off
defparam \Mux49~9 .lut_mask = 16'hBCB0;
defparam \Mux49~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N20
cycloneive_lcell_comb \Mux49~19 (
// Equation(s):
// Mux491 = (instruction_D[18] & ((\Mux49~16_combout  & (\Mux49~18_combout )) # (!\Mux49~16_combout  & ((\Mux49~11_combout ))))) # (!instruction_D[18] & (((\Mux49~16_combout ))))

	.dataa(\Mux49~18_combout ),
	.datab(instruction_D_18),
	.datac(\Mux49~16_combout ),
	.datad(\Mux49~11_combout ),
	.cin(gnd),
	.combout(Mux491),
	.cout());
// synopsys translate_off
defparam \Mux49~19 .lut_mask = 16'hBCB0;
defparam \Mux49~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N14
cycloneive_lcell_comb \Mux50~9 (
// Equation(s):
// Mux50 = (instruction_D[16] & ((\Mux50~6_combout  & ((\Mux50~8_combout ))) # (!\Mux50~6_combout  & (\Mux50~1_combout )))) # (!instruction_D[16] & (\Mux50~6_combout ))

	.dataa(instruction_D_16),
	.datab(\Mux50~6_combout ),
	.datac(\Mux50~1_combout ),
	.datad(\Mux50~8_combout ),
	.cin(gnd),
	.combout(Mux50),
	.cout());
// synopsys translate_off
defparam \Mux50~9 .lut_mask = 16'hEC64;
defparam \Mux50~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N18
cycloneive_lcell_comb \Mux50~19 (
// Equation(s):
// Mux501 = (instruction_D[19] & ((\Mux50~16_combout  & ((\Mux50~18_combout ))) # (!\Mux50~16_combout  & (\Mux50~11_combout )))) # (!instruction_D[19] & (\Mux50~16_combout ))

	.dataa(instruction_D_19),
	.datab(\Mux50~16_combout ),
	.datac(\Mux50~11_combout ),
	.datad(\Mux50~18_combout ),
	.cin(gnd),
	.combout(Mux501),
	.cout());
// synopsys translate_off
defparam \Mux50~19 .lut_mask = 16'hEC64;
defparam \Mux50~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N12
cycloneive_lcell_comb \Mux51~9 (
// Equation(s):
// Mux51 = (instruction_D[16] & ((\Mux51~6_combout  & (\Mux51~8_combout )) # (!\Mux51~6_combout  & ((\Mux51~1_combout ))))) # (!instruction_D[16] & (((\Mux51~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux51~8_combout ),
	.datac(\Mux51~1_combout ),
	.datad(\Mux51~6_combout ),
	.cin(gnd),
	.combout(Mux51),
	.cout());
// synopsys translate_off
defparam \Mux51~9 .lut_mask = 16'hDDA0;
defparam \Mux51~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N10
cycloneive_lcell_comb \Mux51~19 (
// Equation(s):
// Mux511 = (instruction_D[18] & ((\Mux51~16_combout  & (\Mux51~18_combout )) # (!\Mux51~16_combout  & ((\Mux51~11_combout ))))) # (!instruction_D[18] & (((\Mux51~16_combout ))))

	.dataa(instruction_D_18),
	.datab(\Mux51~18_combout ),
	.datac(\Mux51~11_combout ),
	.datad(\Mux51~16_combout ),
	.cin(gnd),
	.combout(Mux511),
	.cout());
// synopsys translate_off
defparam \Mux51~19 .lut_mask = 16'hDDA0;
defparam \Mux51~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N12
cycloneive_lcell_comb \Mux54~9 (
// Equation(s):
// Mux54 = (instruction_D[16] & ((\Mux54~6_combout  & ((\Mux54~8_combout ))) # (!\Mux54~6_combout  & (\Mux54~1_combout )))) # (!instruction_D[16] & (((\Mux54~6_combout ))))

	.dataa(\Mux54~1_combout ),
	.datab(instruction_D_16),
	.datac(\Mux54~8_combout ),
	.datad(\Mux54~6_combout ),
	.cin(gnd),
	.combout(Mux54),
	.cout());
// synopsys translate_off
defparam \Mux54~9 .lut_mask = 16'hF388;
defparam \Mux54~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N4
cycloneive_lcell_comb \Mux54~19 (
// Equation(s):
// Mux541 = (instruction_D[19] & ((\Mux54~16_combout  & (\Mux54~18_combout )) # (!\Mux54~16_combout  & ((\Mux54~11_combout ))))) # (!instruction_D[19] & (((\Mux54~16_combout ))))

	.dataa(\Mux54~18_combout ),
	.datab(instruction_D_19),
	.datac(\Mux54~11_combout ),
	.datad(\Mux54~16_combout ),
	.cin(gnd),
	.combout(Mux541),
	.cout());
// synopsys translate_off
defparam \Mux54~19 .lut_mask = 16'hBBC0;
defparam \Mux54~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N14
cycloneive_lcell_comb \Mux55~9 (
// Equation(s):
// Mux55 = (instruction_D[16] & ((\Mux55~6_combout  & (\Mux55~8_combout )) # (!\Mux55~6_combout  & ((\Mux55~1_combout ))))) # (!instruction_D[16] & (((\Mux55~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux55~8_combout ),
	.datac(\Mux55~6_combout ),
	.datad(\Mux55~1_combout ),
	.cin(gnd),
	.combout(Mux55),
	.cout());
// synopsys translate_off
defparam \Mux55~9 .lut_mask = 16'hDAD0;
defparam \Mux55~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N20
cycloneive_lcell_comb \Mux55~19 (
// Equation(s):
// Mux551 = (instruction_D[18] & ((\Mux55~16_combout  & (\Mux55~18_combout )) # (!\Mux55~16_combout  & ((\Mux55~11_combout ))))) # (!instruction_D[18] & (((\Mux55~16_combout ))))

	.dataa(\Mux55~18_combout ),
	.datab(\Mux55~11_combout ),
	.datac(instruction_D_18),
	.datad(\Mux55~16_combout ),
	.cin(gnd),
	.combout(Mux551),
	.cout());
// synopsys translate_off
defparam \Mux55~19 .lut_mask = 16'hAFC0;
defparam \Mux55~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N24
cycloneive_lcell_comb \Mux52~9 (
// Equation(s):
// Mux52 = (instruction_D[16] & ((\Mux52~6_combout  & (\Mux52~8_combout )) # (!\Mux52~6_combout  & ((\Mux52~1_combout ))))) # (!instruction_D[16] & (((\Mux52~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux52~8_combout ),
	.datac(\Mux52~1_combout ),
	.datad(\Mux52~6_combout ),
	.cin(gnd),
	.combout(Mux52),
	.cout());
// synopsys translate_off
defparam \Mux52~9 .lut_mask = 16'hDDA0;
defparam \Mux52~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N18
cycloneive_lcell_comb \Mux52~19 (
// Equation(s):
// Mux521 = (instruction_D[19] & ((\Mux52~16_combout  & (\Mux52~18_combout )) # (!\Mux52~16_combout  & ((\Mux52~11_combout ))))) # (!instruction_D[19] & (((\Mux52~16_combout ))))

	.dataa(instruction_D_19),
	.datab(\Mux52~18_combout ),
	.datac(\Mux52~16_combout ),
	.datad(\Mux52~11_combout ),
	.cin(gnd),
	.combout(Mux521),
	.cout());
// synopsys translate_off
defparam \Mux52~19 .lut_mask = 16'hDAD0;
defparam \Mux52~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N8
cycloneive_lcell_comb \Mux53~9 (
// Equation(s):
// Mux53 = (instruction_D[16] & ((\Mux53~6_combout  & ((\Mux53~8_combout ))) # (!\Mux53~6_combout  & (\Mux53~1_combout )))) # (!instruction_D[16] & (((\Mux53~6_combout ))))

	.dataa(\Mux53~1_combout ),
	.datab(instruction_D_16),
	.datac(\Mux53~8_combout ),
	.datad(\Mux53~6_combout ),
	.cin(gnd),
	.combout(Mux53),
	.cout());
// synopsys translate_off
defparam \Mux53~9 .lut_mask = 16'hF388;
defparam \Mux53~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N16
cycloneive_lcell_comb \Mux53~19 (
// Equation(s):
// Mux531 = (instruction_D[18] & ((\Mux53~16_combout  & ((\Mux53~18_combout ))) # (!\Mux53~16_combout  & (\Mux53~11_combout )))) # (!instruction_D[18] & (((\Mux53~16_combout ))))

	.dataa(instruction_D_18),
	.datab(\Mux53~11_combout ),
	.datac(\Mux53~18_combout ),
	.datad(\Mux53~16_combout ),
	.cin(gnd),
	.combout(Mux531),
	.cout());
// synopsys translate_off
defparam \Mux53~19 .lut_mask = 16'hF588;
defparam \Mux53~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N16
cycloneive_lcell_comb \Mux56~9 (
// Equation(s):
// Mux56 = (instruction_D[16] & ((\Mux56~6_combout  & ((\Mux56~8_combout ))) # (!\Mux56~6_combout  & (\Mux56~1_combout )))) # (!instruction_D[16] & (((\Mux56~6_combout ))))

	.dataa(\Mux56~1_combout ),
	.datab(instruction_D_16),
	.datac(\Mux56~8_combout ),
	.datad(\Mux56~6_combout ),
	.cin(gnd),
	.combout(Mux56),
	.cout());
// synopsys translate_off
defparam \Mux56~9 .lut_mask = 16'hF388;
defparam \Mux56~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N4
cycloneive_lcell_comb \Mux56~19 (
// Equation(s):
// Mux561 = (instruction_D[19] & ((\Mux56~16_combout  & (\Mux56~18_combout )) # (!\Mux56~16_combout  & ((\Mux56~11_combout ))))) # (!instruction_D[19] & (((\Mux56~16_combout ))))

	.dataa(\Mux56~18_combout ),
	.datab(instruction_D_19),
	.datac(\Mux56~16_combout ),
	.datad(\Mux56~11_combout ),
	.cin(gnd),
	.combout(Mux561),
	.cout());
// synopsys translate_off
defparam \Mux56~19 .lut_mask = 16'hBCB0;
defparam \Mux56~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N26
cycloneive_lcell_comb \Mux57~9 (
// Equation(s):
// Mux57 = (instruction_D[16] & ((\Mux57~6_combout  & ((\Mux57~8_combout ))) # (!\Mux57~6_combout  & (\Mux57~1_combout )))) # (!instruction_D[16] & (((\Mux57~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux57~1_combout ),
	.datac(\Mux57~6_combout ),
	.datad(\Mux57~8_combout ),
	.cin(gnd),
	.combout(Mux57),
	.cout());
// synopsys translate_off
defparam \Mux57~9 .lut_mask = 16'hF858;
defparam \Mux57~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N2
cycloneive_lcell_comb \Mux57~19 (
// Equation(s):
// Mux571 = (instruction_D[18] & ((\Mux57~16_combout  & ((\Mux57~18_combout ))) # (!\Mux57~16_combout  & (\Mux57~11_combout )))) # (!instruction_D[18] & (((\Mux57~16_combout ))))

	.dataa(\Mux57~11_combout ),
	.datab(\Mux57~18_combout ),
	.datac(instruction_D_18),
	.datad(\Mux57~16_combout ),
	.cin(gnd),
	.combout(Mux571),
	.cout());
// synopsys translate_off
defparam \Mux57~19 .lut_mask = 16'hCFA0;
defparam \Mux57~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N20
cycloneive_lcell_comb \Mux58~9 (
// Equation(s):
// Mux58 = (instruction_D[16] & ((\Mux58~6_combout  & (\Mux58~8_combout )) # (!\Mux58~6_combout  & ((\Mux58~1_combout ))))) # (!instruction_D[16] & (((\Mux58~6_combout ))))

	.dataa(\Mux58~8_combout ),
	.datab(instruction_D_16),
	.datac(\Mux58~1_combout ),
	.datad(\Mux58~6_combout ),
	.cin(gnd),
	.combout(Mux58),
	.cout());
// synopsys translate_off
defparam \Mux58~9 .lut_mask = 16'hBBC0;
defparam \Mux58~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N10
cycloneive_lcell_comb \Mux58~19 (
// Equation(s):
// Mux581 = (instruction_D[19] & ((\Mux58~16_combout  & ((\Mux58~18_combout ))) # (!\Mux58~16_combout  & (\Mux58~11_combout )))) # (!instruction_D[19] & (((\Mux58~16_combout ))))

	.dataa(\Mux58~11_combout ),
	.datab(instruction_D_19),
	.datac(\Mux58~18_combout ),
	.datad(\Mux58~16_combout ),
	.cin(gnd),
	.combout(Mux581),
	.cout());
// synopsys translate_off
defparam \Mux58~19 .lut_mask = 16'hF388;
defparam \Mux58~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N6
cycloneive_lcell_comb \Mux29~9 (
// Equation(s):
// Mux29 = (instruction_D[21] & ((\Mux29~6_combout  & ((\Mux29~8_combout ))) # (!\Mux29~6_combout  & (\Mux29~1_combout )))) # (!instruction_D[21] & (((\Mux29~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux29~1_combout ),
	.datac(\Mux29~8_combout ),
	.datad(\Mux29~6_combout ),
	.cin(gnd),
	.combout(Mux29),
	.cout());
// synopsys translate_off
defparam \Mux29~9 .lut_mask = 16'hF588;
defparam \Mux29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N16
cycloneive_lcell_comb \Mux29~19 (
// Equation(s):
// Mux291 = (instruction_D[24] & ((\Mux29~16_combout  & ((\Mux29~18_combout ))) # (!\Mux29~16_combout  & (\Mux29~11_combout )))) # (!instruction_D[24] & (((\Mux29~16_combout ))))

	.dataa(\Mux29~11_combout ),
	.datab(instruction_D_24),
	.datac(\Mux29~18_combout ),
	.datad(\Mux29~16_combout ),
	.cin(gnd),
	.combout(Mux291),
	.cout());
// synopsys translate_off
defparam \Mux29~19 .lut_mask = 16'hF388;
defparam \Mux29~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N26
cycloneive_lcell_comb \Mux30~9 (
// Equation(s):
// Mux30 = (instruction_D[21] & ((\Mux30~6_combout  & (\Mux30~8_combout )) # (!\Mux30~6_combout  & ((\Mux30~1_combout ))))) # (!instruction_D[21] & (\Mux30~6_combout ))

	.dataa(instruction_D_21),
	.datab(\Mux30~6_combout ),
	.datac(\Mux30~8_combout ),
	.datad(\Mux30~1_combout ),
	.cin(gnd),
	.combout(Mux30),
	.cout());
// synopsys translate_off
defparam \Mux30~9 .lut_mask = 16'hE6C4;
defparam \Mux30~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N0
cycloneive_lcell_comb \Mux30~19 (
// Equation(s):
// Mux301 = (instruction_D[24] & ((\Mux30~16_combout  & ((\Mux30~18_combout ))) # (!\Mux30~16_combout  & (\Mux30~11_combout )))) # (!instruction_D[24] & (((\Mux30~16_combout ))))

	.dataa(instruction_D_24),
	.datab(\Mux30~11_combout ),
	.datac(\Mux30~18_combout ),
	.datad(\Mux30~16_combout ),
	.cin(gnd),
	.combout(Mux301),
	.cout());
// synopsys translate_off
defparam \Mux30~19 .lut_mask = 16'hF588;
defparam \Mux30~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N30
cycloneive_lcell_comb \Mux63~9 (
// Equation(s):
// Mux63 = (instruction_D[16] & ((\Mux63~6_combout  & ((\Mux63~8_combout ))) # (!\Mux63~6_combout  & (\Mux63~1_combout )))) # (!instruction_D[16] & (((\Mux63~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux63~1_combout ),
	.datac(\Mux63~8_combout ),
	.datad(\Mux63~6_combout ),
	.cin(gnd),
	.combout(Mux63),
	.cout());
// synopsys translate_off
defparam \Mux63~9 .lut_mask = 16'hF588;
defparam \Mux63~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N10
cycloneive_lcell_comb \Mux63~19 (
// Equation(s):
// Mux631 = (\Mux63~16_combout  & (((\Mux63~18_combout )) # (!instruction_D[18]))) # (!\Mux63~16_combout  & (instruction_D[18] & ((\Mux63~11_combout ))))

	.dataa(\Mux63~16_combout ),
	.datab(instruction_D_18),
	.datac(\Mux63~18_combout ),
	.datad(\Mux63~11_combout ),
	.cin(gnd),
	.combout(Mux631),
	.cout());
// synopsys translate_off
defparam \Mux63~19 .lut_mask = 16'hE6A2;
defparam \Mux63~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N2
cycloneive_lcell_comb \Mux62~9 (
// Equation(s):
// Mux62 = (instruction_D[16] & ((\Mux62~6_combout  & ((\Mux62~8_combout ))) # (!\Mux62~6_combout  & (\Mux62~1_combout )))) # (!instruction_D[16] & (((\Mux62~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux62~1_combout ),
	.datac(\Mux62~6_combout ),
	.datad(\Mux62~8_combout ),
	.cin(gnd),
	.combout(Mux62),
	.cout());
// synopsys translate_off
defparam \Mux62~9 .lut_mask = 16'hF858;
defparam \Mux62~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N22
cycloneive_lcell_comb \Mux62~19 (
// Equation(s):
// Mux621 = (instruction_D[19] & ((\Mux62~16_combout  & ((\Mux62~18_combout ))) # (!\Mux62~16_combout  & (\Mux62~11_combout )))) # (!instruction_D[19] & (((\Mux62~16_combout ))))

	.dataa(instruction_D_19),
	.datab(\Mux62~11_combout ),
	.datac(\Mux62~18_combout ),
	.datad(\Mux62~16_combout ),
	.cin(gnd),
	.combout(Mux621),
	.cout());
// synopsys translate_off
defparam \Mux62~19 .lut_mask = 16'hF588;
defparam \Mux62~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N20
cycloneive_lcell_comb \Mux27~9 (
// Equation(s):
// Mux27 = (instruction_D[21] & ((\Mux27~6_combout  & (\Mux27~8_combout )) # (!\Mux27~6_combout  & ((\Mux27~1_combout ))))) # (!instruction_D[21] & (((\Mux27~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux27~8_combout ),
	.datac(\Mux27~1_combout ),
	.datad(\Mux27~6_combout ),
	.cin(gnd),
	.combout(Mux27),
	.cout());
// synopsys translate_off
defparam \Mux27~9 .lut_mask = 16'hDDA0;
defparam \Mux27~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N22
cycloneive_lcell_comb \Mux27~19 (
// Equation(s):
// Mux271 = (instruction_D[23] & ((\Mux27~16_combout  & (\Mux27~18_combout )) # (!\Mux27~16_combout  & ((\Mux27~11_combout ))))) # (!instruction_D[23] & (((\Mux27~16_combout ))))

	.dataa(instruction_D_23),
	.datab(\Mux27~18_combout ),
	.datac(\Mux27~11_combout ),
	.datad(\Mux27~16_combout ),
	.cin(gnd),
	.combout(Mux271),
	.cout());
// synopsys translate_off
defparam \Mux27~19 .lut_mask = 16'hDDA0;
defparam \Mux27~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N30
cycloneive_lcell_comb \Mux28~9 (
// Equation(s):
// Mux28 = (instruction_D[21] & ((\Mux28~6_combout  & (\Mux28~8_combout )) # (!\Mux28~6_combout  & ((\Mux28~1_combout ))))) # (!instruction_D[21] & (((\Mux28~6_combout ))))

	.dataa(\Mux28~8_combout ),
	.datab(instruction_D_21),
	.datac(\Mux28~1_combout ),
	.datad(\Mux28~6_combout ),
	.cin(gnd),
	.combout(Mux28),
	.cout());
// synopsys translate_off
defparam \Mux28~9 .lut_mask = 16'hBBC0;
defparam \Mux28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N24
cycloneive_lcell_comb \Mux28~19 (
// Equation(s):
// Mux281 = (instruction_D[23] & ((\Mux28~16_combout  & (\Mux28~18_combout )) # (!\Mux28~16_combout  & ((\Mux28~11_combout ))))) # (!instruction_D[23] & (((\Mux28~16_combout ))))

	.dataa(instruction_D_23),
	.datab(\Mux28~18_combout ),
	.datac(\Mux28~11_combout ),
	.datad(\Mux28~16_combout ),
	.cin(gnd),
	.combout(Mux281),
	.cout());
// synopsys translate_off
defparam \Mux28~19 .lut_mask = 16'hDDA0;
defparam \Mux28~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N30
cycloneive_lcell_comb \Mux61~9 (
// Equation(s):
// Mux61 = (instruction_D[16] & ((\Mux61~6_combout  & ((\Mux61~8_combout ))) # (!\Mux61~6_combout  & (\Mux61~1_combout )))) # (!instruction_D[16] & (((\Mux61~6_combout ))))

	.dataa(\Mux61~1_combout ),
	.datab(instruction_D_16),
	.datac(\Mux61~8_combout ),
	.datad(\Mux61~6_combout ),
	.cin(gnd),
	.combout(Mux61),
	.cout());
// synopsys translate_off
defparam \Mux61~9 .lut_mask = 16'hF388;
defparam \Mux61~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N12
cycloneive_lcell_comb \Mux61~19 (
// Equation(s):
// Mux611 = (\Mux61~16_combout  & (((\Mux61~18_combout )) # (!instruction_D[18]))) # (!\Mux61~16_combout  & (instruction_D[18] & (\Mux61~11_combout )))

	.dataa(\Mux61~16_combout ),
	.datab(instruction_D_18),
	.datac(\Mux61~11_combout ),
	.datad(\Mux61~18_combout ),
	.cin(gnd),
	.combout(Mux611),
	.cout());
// synopsys translate_off
defparam \Mux61~19 .lut_mask = 16'hEA62;
defparam \Mux61~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N26
cycloneive_lcell_comb \Mux23~9 (
// Equation(s):
// Mux23 = (instruction_D[21] & ((\Mux23~6_combout  & ((\Mux23~8_combout ))) # (!\Mux23~6_combout  & (\Mux23~1_combout )))) # (!instruction_D[21] & (((\Mux23~6_combout ))))

	.dataa(\Mux23~1_combout ),
	.datab(instruction_D_21),
	.datac(\Mux23~8_combout ),
	.datad(\Mux23~6_combout ),
	.cin(gnd),
	.combout(Mux23),
	.cout());
// synopsys translate_off
defparam \Mux23~9 .lut_mask = 16'hF388;
defparam \Mux23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N26
cycloneive_lcell_comb \Mux23~19 (
// Equation(s):
// Mux231 = (instruction_D[23] & ((\Mux23~16_combout  & ((\Mux23~18_combout ))) # (!\Mux23~16_combout  & (\Mux23~11_combout )))) # (!instruction_D[23] & (((\Mux23~16_combout ))))

	.dataa(instruction_D_23),
	.datab(\Mux23~11_combout ),
	.datac(\Mux23~16_combout ),
	.datad(\Mux23~18_combout ),
	.cin(gnd),
	.combout(Mux231),
	.cout());
// synopsys translate_off
defparam \Mux23~19 .lut_mask = 16'hF858;
defparam \Mux23~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N20
cycloneive_lcell_comb \Mux24~9 (
// Equation(s):
// Mux24 = (instruction_D[21] & ((\Mux24~6_combout  & ((\Mux24~8_combout ))) # (!\Mux24~6_combout  & (\Mux24~1_combout )))) # (!instruction_D[21] & (((\Mux24~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux24~1_combout ),
	.datac(\Mux24~8_combout ),
	.datad(\Mux24~6_combout ),
	.cin(gnd),
	.combout(Mux24),
	.cout());
// synopsys translate_off
defparam \Mux24~9 .lut_mask = 16'hF588;
defparam \Mux24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N4
cycloneive_lcell_comb \Mux24~19 (
// Equation(s):
// Mux241 = (instruction_D[24] & ((\Mux24~16_combout  & (\Mux24~18_combout )) # (!\Mux24~16_combout  & ((\Mux24~11_combout ))))) # (!instruction_D[24] & (((\Mux24~16_combout ))))

	.dataa(\Mux24~18_combout ),
	.datab(\Mux24~11_combout ),
	.datac(instruction_D_24),
	.datad(\Mux24~16_combout ),
	.cin(gnd),
	.combout(Mux241),
	.cout());
// synopsys translate_off
defparam \Mux24~19 .lut_mask = 16'hAFC0;
defparam \Mux24~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N14
cycloneive_lcell_comb \Mux25~9 (
// Equation(s):
// Mux25 = (instruction_D[21] & ((\Mux25~6_combout  & ((\Mux25~8_combout ))) # (!\Mux25~6_combout  & (\Mux25~1_combout )))) # (!instruction_D[21] & (((\Mux25~6_combout ))))

	.dataa(\Mux25~1_combout ),
	.datab(instruction_D_21),
	.datac(\Mux25~8_combout ),
	.datad(\Mux25~6_combout ),
	.cin(gnd),
	.combout(Mux25),
	.cout());
// synopsys translate_off
defparam \Mux25~9 .lut_mask = 16'hF388;
defparam \Mux25~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N18
cycloneive_lcell_comb \Mux25~19 (
// Equation(s):
// Mux251 = (instruction_D[23] & ((\Mux25~16_combout  & ((\Mux25~18_combout ))) # (!\Mux25~16_combout  & (\Mux25~11_combout )))) # (!instruction_D[23] & (((\Mux25~16_combout ))))

	.dataa(instruction_D_23),
	.datab(\Mux25~11_combout ),
	.datac(\Mux25~16_combout ),
	.datad(\Mux25~18_combout ),
	.cin(gnd),
	.combout(Mux251),
	.cout());
// synopsys translate_off
defparam \Mux25~19 .lut_mask = 16'hF858;
defparam \Mux25~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N10
cycloneive_lcell_comb \Mux26~9 (
// Equation(s):
// Mux26 = (instruction_D[21] & ((\Mux26~6_combout  & (\Mux26~8_combout )) # (!\Mux26~6_combout  & ((\Mux26~1_combout ))))) # (!instruction_D[21] & (((\Mux26~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux26~8_combout ),
	.datac(\Mux26~6_combout ),
	.datad(\Mux26~1_combout ),
	.cin(gnd),
	.combout(Mux26),
	.cout());
// synopsys translate_off
defparam \Mux26~9 .lut_mask = 16'hDAD0;
defparam \Mux26~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N28
cycloneive_lcell_comb \Mux26~19 (
// Equation(s):
// Mux261 = (\Mux26~16_combout  & (((\Mux26~18_combout )) # (!instruction_D[24]))) # (!\Mux26~16_combout  & (instruction_D[24] & (\Mux26~11_combout )))

	.dataa(\Mux26~16_combout ),
	.datab(instruction_D_24),
	.datac(\Mux26~11_combout ),
	.datad(\Mux26~18_combout ),
	.cin(gnd),
	.combout(Mux261),
	.cout());
// synopsys translate_off
defparam \Mux26~19 .lut_mask = 16'hEA62;
defparam \Mux26~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N14
cycloneive_lcell_comb \Mux60~9 (
// Equation(s):
// Mux60 = (instruction_D[16] & ((\Mux60~6_combout  & (\Mux60~8_combout )) # (!\Mux60~6_combout  & ((\Mux60~1_combout ))))) # (!instruction_D[16] & (((\Mux60~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux60~8_combout ),
	.datac(\Mux60~1_combout ),
	.datad(\Mux60~6_combout ),
	.cin(gnd),
	.combout(Mux60),
	.cout());
// synopsys translate_off
defparam \Mux60~9 .lut_mask = 16'hDDA0;
defparam \Mux60~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N20
cycloneive_lcell_comb \Mux60~19 (
// Equation(s):
// Mux601 = (\Mux60~16_combout  & (((\Mux60~18_combout )) # (!instruction_D[19]))) # (!\Mux60~16_combout  & (instruction_D[19] & (\Mux60~11_combout )))

	.dataa(\Mux60~16_combout ),
	.datab(instruction_D_19),
	.datac(\Mux60~11_combout ),
	.datad(\Mux60~18_combout ),
	.cin(gnd),
	.combout(Mux601),
	.cout());
// synopsys translate_off
defparam \Mux60~19 .lut_mask = 16'hEA62;
defparam \Mux60~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N4
cycloneive_lcell_comb \Mux15~9 (
// Equation(s):
// Mux15 = (instruction_D[21] & ((\Mux15~6_combout  & (\Mux15~8_combout )) # (!\Mux15~6_combout  & ((\Mux15~1_combout ))))) # (!instruction_D[21] & (((\Mux15~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux15~8_combout ),
	.datac(\Mux15~6_combout ),
	.datad(\Mux15~1_combout ),
	.cin(gnd),
	.combout(Mux15),
	.cout());
// synopsys translate_off
defparam \Mux15~9 .lut_mask = 16'hDAD0;
defparam \Mux15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N12
cycloneive_lcell_comb \Mux15~19 (
// Equation(s):
// Mux151 = (instruction_D[23] & ((\Mux15~16_combout  & ((\Mux15~18_combout ))) # (!\Mux15~16_combout  & (\Mux15~11_combout )))) # (!instruction_D[23] & (((\Mux15~16_combout ))))

	.dataa(\Mux15~11_combout ),
	.datab(instruction_D_23),
	.datac(\Mux15~16_combout ),
	.datad(\Mux15~18_combout ),
	.cin(gnd),
	.combout(Mux151),
	.cout());
// synopsys translate_off
defparam \Mux15~19 .lut_mask = 16'hF838;
defparam \Mux15~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N8
cycloneive_lcell_comb \Mux16~9 (
// Equation(s):
// Mux16 = (instruction_D[21] & ((\Mux16~6_combout  & (\Mux16~8_combout )) # (!\Mux16~6_combout  & ((\Mux16~1_combout ))))) # (!instruction_D[21] & (((\Mux16~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux16~8_combout ),
	.datac(\Mux16~1_combout ),
	.datad(\Mux16~6_combout ),
	.cin(gnd),
	.combout(Mux16),
	.cout());
// synopsys translate_off
defparam \Mux16~9 .lut_mask = 16'hDDA0;
defparam \Mux16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N16
cycloneive_lcell_comb \Mux16~19 (
// Equation(s):
// Mux161 = (instruction_D[24] & ((\Mux16~16_combout  & (\Mux16~18_combout )) # (!\Mux16~16_combout  & ((\Mux16~11_combout ))))) # (!instruction_D[24] & (((\Mux16~16_combout ))))

	.dataa(\Mux16~18_combout ),
	.datab(instruction_D_24),
	.datac(\Mux16~11_combout ),
	.datad(\Mux16~16_combout ),
	.cin(gnd),
	.combout(Mux161),
	.cout());
// synopsys translate_off
defparam \Mux16~19 .lut_mask = 16'hBBC0;
defparam \Mux16~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N12
cycloneive_lcell_comb \Mux17~9 (
// Equation(s):
// Mux17 = (instruction_D[21] & ((\Mux17~6_combout  & (\Mux17~8_combout )) # (!\Mux17~6_combout  & ((\Mux17~1_combout ))))) # (!instruction_D[21] & (((\Mux17~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux17~8_combout ),
	.datac(\Mux17~6_combout ),
	.datad(\Mux17~1_combout ),
	.cin(gnd),
	.combout(Mux17),
	.cout());
// synopsys translate_off
defparam \Mux17~9 .lut_mask = 16'hDAD0;
defparam \Mux17~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N20
cycloneive_lcell_comb \Mux17~19 (
// Equation(s):
// Mux171 = (instruction_D[23] & ((\Mux17~16_combout  & ((\Mux17~18_combout ))) # (!\Mux17~16_combout  & (\Mux17~11_combout )))) # (!instruction_D[23] & (((\Mux17~16_combout ))))

	.dataa(instruction_D_23),
	.datab(\Mux17~11_combout ),
	.datac(\Mux17~18_combout ),
	.datad(\Mux17~16_combout ),
	.cin(gnd),
	.combout(Mux171),
	.cout());
// synopsys translate_off
defparam \Mux17~19 .lut_mask = 16'hF588;
defparam \Mux17~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N10
cycloneive_lcell_comb \Mux18~9 (
// Equation(s):
// Mux18 = (instruction_D[21] & ((\Mux18~6_combout  & (\Mux18~8_combout )) # (!\Mux18~6_combout  & ((\Mux18~1_combout ))))) # (!instruction_D[21] & (((\Mux18~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux18~8_combout ),
	.datac(\Mux18~1_combout ),
	.datad(\Mux18~6_combout ),
	.cin(gnd),
	.combout(Mux18),
	.cout());
// synopsys translate_off
defparam \Mux18~9 .lut_mask = 16'hDDA0;
defparam \Mux18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N10
cycloneive_lcell_comb \Mux18~19 (
// Equation(s):
// Mux181 = (\Mux18~16_combout  & ((\Mux18~18_combout ) # ((!instruction_D[24])))) # (!\Mux18~16_combout  & (((instruction_D[24] & \Mux18~11_combout ))))

	.dataa(\Mux18~18_combout ),
	.datab(\Mux18~16_combout ),
	.datac(instruction_D_24),
	.datad(\Mux18~11_combout ),
	.cin(gnd),
	.combout(Mux181),
	.cout());
// synopsys translate_off
defparam \Mux18~19 .lut_mask = 16'hBC8C;
defparam \Mux18~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N24
cycloneive_lcell_comb \Mux19~9 (
// Equation(s):
// Mux19 = (instruction_D[21] & ((\Mux19~6_combout  & (\Mux19~8_combout )) # (!\Mux19~6_combout  & ((\Mux19~1_combout ))))) # (!instruction_D[21] & (((\Mux19~6_combout ))))

	.dataa(\Mux19~8_combout ),
	.datab(instruction_D_21),
	.datac(\Mux19~1_combout ),
	.datad(\Mux19~6_combout ),
	.cin(gnd),
	.combout(Mux19),
	.cout());
// synopsys translate_off
defparam \Mux19~9 .lut_mask = 16'hBBC0;
defparam \Mux19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N22
cycloneive_lcell_comb \Mux19~19 (
// Equation(s):
// Mux191 = (instruction_D[23] & ((\Mux19~16_combout  & ((\Mux19~18_combout ))) # (!\Mux19~16_combout  & (\Mux19~11_combout )))) # (!instruction_D[23] & (((\Mux19~16_combout ))))

	.dataa(instruction_D_23),
	.datab(\Mux19~11_combout ),
	.datac(\Mux19~16_combout ),
	.datad(\Mux19~18_combout ),
	.cin(gnd),
	.combout(Mux191),
	.cout());
// synopsys translate_off
defparam \Mux19~19 .lut_mask = 16'hF858;
defparam \Mux19~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N6
cycloneive_lcell_comb \Mux20~9 (
// Equation(s):
// Mux20 = (instruction_D[21] & ((\Mux20~6_combout  & ((\Mux20~8_combout ))) # (!\Mux20~6_combout  & (\Mux20~1_combout )))) # (!instruction_D[21] & (((\Mux20~6_combout ))))

	.dataa(\Mux20~1_combout ),
	.datab(instruction_D_21),
	.datac(\Mux20~8_combout ),
	.datad(\Mux20~6_combout ),
	.cin(gnd),
	.combout(Mux20),
	.cout());
// synopsys translate_off
defparam \Mux20~9 .lut_mask = 16'hF388;
defparam \Mux20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N4
cycloneive_lcell_comb \Mux20~19 (
// Equation(s):
// Mux201 = (\Mux20~16_combout  & ((\Mux20~18_combout ) # ((!instruction_D[24])))) # (!\Mux20~16_combout  & (((instruction_D[24] & \Mux20~11_combout ))))

	.dataa(\Mux20~18_combout ),
	.datab(\Mux20~16_combout ),
	.datac(instruction_D_24),
	.datad(\Mux20~11_combout ),
	.cin(gnd),
	.combout(Mux201),
	.cout());
// synopsys translate_off
defparam \Mux20~19 .lut_mask = 16'hBC8C;
defparam \Mux20~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N12
cycloneive_lcell_comb \Mux21~9 (
// Equation(s):
// Mux21 = (instruction_D[21] & ((\Mux21~6_combout  & ((\Mux21~8_combout ))) # (!\Mux21~6_combout  & (\Mux21~1_combout )))) # (!instruction_D[21] & (((\Mux21~6_combout ))))

	.dataa(\Mux21~1_combout ),
	.datab(\Mux21~8_combout ),
	.datac(instruction_D_21),
	.datad(\Mux21~6_combout ),
	.cin(gnd),
	.combout(Mux21),
	.cout());
// synopsys translate_off
defparam \Mux21~9 .lut_mask = 16'hCFA0;
defparam \Mux21~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N8
cycloneive_lcell_comb \Mux21~19 (
// Equation(s):
// Mux211 = (instruction_D[23] & ((\Mux21~16_combout  & ((\Mux21~18_combout ))) # (!\Mux21~16_combout  & (\Mux21~11_combout )))) # (!instruction_D[23] & (((\Mux21~16_combout ))))

	.dataa(\Mux21~11_combout ),
	.datab(\Mux21~18_combout ),
	.datac(instruction_D_23),
	.datad(\Mux21~16_combout ),
	.cin(gnd),
	.combout(Mux211),
	.cout());
// synopsys translate_off
defparam \Mux21~19 .lut_mask = 16'hCFA0;
defparam \Mux21~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N22
cycloneive_lcell_comb \Mux22~9 (
// Equation(s):
// Mux22 = (\Mux22~6_combout  & (((\Mux22~8_combout )) # (!instruction_D[21]))) # (!\Mux22~6_combout  & (instruction_D[21] & ((\Mux22~1_combout ))))

	.dataa(\Mux22~6_combout ),
	.datab(instruction_D_21),
	.datac(\Mux22~8_combout ),
	.datad(\Mux22~1_combout ),
	.cin(gnd),
	.combout(Mux22),
	.cout());
// synopsys translate_off
defparam \Mux22~9 .lut_mask = 16'hE6A2;
defparam \Mux22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N22
cycloneive_lcell_comb \Mux22~19 (
// Equation(s):
// Mux221 = (instruction_D[24] & ((\Mux22~16_combout  & ((\Mux22~18_combout ))) # (!\Mux22~16_combout  & (\Mux22~11_combout )))) # (!instruction_D[24] & (((\Mux22~16_combout ))))

	.dataa(instruction_D_24),
	.datab(\Mux22~11_combout ),
	.datac(\Mux22~16_combout ),
	.datad(\Mux22~18_combout ),
	.cin(gnd),
	.combout(Mux221),
	.cout());
// synopsys translate_off
defparam \Mux22~19 .lut_mask = 16'hF858;
defparam \Mux22~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N24
cycloneive_lcell_comb \Mux59~9 (
// Equation(s):
// Mux59 = (instruction_D[16] & ((\Mux59~6_combout  & (\Mux59~8_combout )) # (!\Mux59~6_combout  & ((\Mux59~1_combout ))))) # (!instruction_D[16] & (((\Mux59~6_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux59~8_combout ),
	.datac(\Mux59~1_combout ),
	.datad(\Mux59~6_combout ),
	.cin(gnd),
	.combout(Mux59),
	.cout());
// synopsys translate_off
defparam \Mux59~9 .lut_mask = 16'hDDA0;
defparam \Mux59~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N14
cycloneive_lcell_comb \Mux59~19 (
// Equation(s):
// Mux591 = (instruction_D[18] & ((\Mux59~16_combout  & (\Mux59~18_combout )) # (!\Mux59~16_combout  & ((\Mux59~11_combout ))))) # (!instruction_D[18] & (((\Mux59~16_combout ))))

	.dataa(instruction_D_18),
	.datab(\Mux59~18_combout ),
	.datac(\Mux59~16_combout ),
	.datad(\Mux59~11_combout ),
	.cin(gnd),
	.combout(Mux591),
	.cout());
// synopsys translate_off
defparam \Mux59~19 .lut_mask = 16'hDAD0;
defparam \Mux59~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N8
cycloneive_lcell_comb \Mux0~9 (
// Equation(s):
// Mux0 = (instruction_D[21] & ((\Mux0~6_combout  & ((\Mux0~8_combout ))) # (!\Mux0~6_combout  & (\Mux0~1_combout )))) # (!instruction_D[21] & (((\Mux0~6_combout ))))

	.dataa(\Mux0~1_combout ),
	.datab(instruction_D_21),
	.datac(\Mux0~6_combout ),
	.datad(\Mux0~8_combout ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
// synopsys translate_off
defparam \Mux0~9 .lut_mask = 16'hF838;
defparam \Mux0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N4
cycloneive_lcell_comb \Mux0~19 (
// Equation(s):
// Mux01 = (instruction_D[24] & ((\Mux0~16_combout  & ((\Mux0~18_combout ))) # (!\Mux0~16_combout  & (\Mux0~11_combout )))) # (!instruction_D[24] & (((\Mux0~16_combout ))))

	.dataa(instruction_D_24),
	.datab(\Mux0~11_combout ),
	.datac(\Mux0~18_combout ),
	.datad(\Mux0~16_combout ),
	.cin(gnd),
	.combout(Mux01),
	.cout());
// synopsys translate_off
defparam \Mux0~19 .lut_mask = 16'hF588;
defparam \Mux0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N6
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// Mux2 = (instruction_D[21] & ((\Mux2~6_combout  & (\Mux2~8_combout )) # (!\Mux2~6_combout  & ((\Mux2~1_combout ))))) # (!instruction_D[21] & (((\Mux2~6_combout ))))

	.dataa(\Mux2~8_combout ),
	.datab(instruction_D_21),
	.datac(\Mux2~1_combout ),
	.datad(\Mux2~6_combout ),
	.cin(gnd),
	.combout(Mux2),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'hBBC0;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N6
cycloneive_lcell_comb \Mux2~19 (
// Equation(s):
// Mux210 = (instruction_D[24] & ((\Mux2~16_combout  & (\Mux2~18_combout )) # (!\Mux2~16_combout  & ((\Mux2~11_combout ))))) # (!instruction_D[24] & (((\Mux2~16_combout ))))

	.dataa(instruction_D_24),
	.datab(\Mux2~18_combout ),
	.datac(\Mux2~11_combout ),
	.datad(\Mux2~16_combout ),
	.cin(gnd),
	.combout(Mux210),
	.cout());
// synopsys translate_off
defparam \Mux2~19 .lut_mask = 16'hDDA0;
defparam \Mux2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N22
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// Mux1 = (\Mux1~6_combout  & (((\Mux1~8_combout )) # (!instruction_D[21]))) # (!\Mux1~6_combout  & (instruction_D[21] & ((\Mux1~1_combout ))))

	.dataa(\Mux1~6_combout ),
	.datab(instruction_D_21),
	.datac(\Mux1~8_combout ),
	.datad(\Mux1~1_combout ),
	.cin(gnd),
	.combout(Mux1),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'hE6A2;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N0
cycloneive_lcell_comb \Mux1~19 (
// Equation(s):
// Mux11 = (instruction_D[23] & ((\Mux1~16_combout  & (\Mux1~18_combout )) # (!\Mux1~16_combout  & ((\Mux1~11_combout ))))) # (!instruction_D[23] & (((\Mux1~16_combout ))))

	.dataa(instruction_D_23),
	.datab(\Mux1~18_combout ),
	.datac(\Mux1~11_combout ),
	.datad(\Mux1~16_combout ),
	.cin(gnd),
	.combout(Mux11),
	.cout());
// synopsys translate_off
defparam \Mux1~19 .lut_mask = 16'hDDA0;
defparam \Mux1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N4
cycloneive_lcell_comb \Mux3~9 (
// Equation(s):
// Mux3 = (instruction_D[21] & ((\Mux3~6_combout  & ((\Mux3~8_combout ))) # (!\Mux3~6_combout  & (\Mux3~1_combout )))) # (!instruction_D[21] & (((\Mux3~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux3~1_combout ),
	.datac(\Mux3~8_combout ),
	.datad(\Mux3~6_combout ),
	.cin(gnd),
	.combout(Mux3),
	.cout());
// synopsys translate_off
defparam \Mux3~9 .lut_mask = 16'hF588;
defparam \Mux3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N12
cycloneive_lcell_comb \Mux3~19 (
// Equation(s):
// Mux31 = (instruction_D[23] & ((\Mux3~16_combout  & ((\Mux3~18_combout ))) # (!\Mux3~16_combout  & (\Mux3~11_combout )))) # (!instruction_D[23] & (((\Mux3~16_combout ))))

	.dataa(\Mux3~11_combout ),
	.datab(instruction_D_23),
	.datac(\Mux3~18_combout ),
	.datad(\Mux3~16_combout ),
	.cin(gnd),
	.combout(Mux31),
	.cout());
// synopsys translate_off
defparam \Mux3~19 .lut_mask = 16'hF388;
defparam \Mux3~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N14
cycloneive_lcell_comb \Mux4~9 (
// Equation(s):
// Mux4 = (instruction_D[21] & ((\Mux4~6_combout  & ((\Mux4~8_combout ))) # (!\Mux4~6_combout  & (\Mux4~1_combout )))) # (!instruction_D[21] & (((\Mux4~6_combout ))))

	.dataa(\Mux4~1_combout ),
	.datab(instruction_D_21),
	.datac(\Mux4~8_combout ),
	.datad(\Mux4~6_combout ),
	.cin(gnd),
	.combout(Mux4),
	.cout());
// synopsys translate_off
defparam \Mux4~9 .lut_mask = 16'hF388;
defparam \Mux4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N2
cycloneive_lcell_comb \Mux4~19 (
// Equation(s):
// Mux410 = (instruction_D[24] & ((\Mux4~16_combout  & (\Mux4~18_combout )) # (!\Mux4~16_combout  & ((\Mux4~11_combout ))))) # (!instruction_D[24] & (((\Mux4~16_combout ))))

	.dataa(\Mux4~18_combout ),
	.datab(instruction_D_24),
	.datac(\Mux4~11_combout ),
	.datad(\Mux4~16_combout ),
	.cin(gnd),
	.combout(Mux410),
	.cout());
// synopsys translate_off
defparam \Mux4~19 .lut_mask = 16'hBBC0;
defparam \Mux4~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N4
cycloneive_lcell_comb \Mux5~9 (
// Equation(s):
// Mux5 = (instruction_D[21] & ((\Mux5~6_combout  & ((\Mux5~8_combout ))) # (!\Mux5~6_combout  & (\Mux5~1_combout )))) # (!instruction_D[21] & (((\Mux5~6_combout ))))

	.dataa(\Mux5~1_combout ),
	.datab(instruction_D_21),
	.datac(\Mux5~8_combout ),
	.datad(\Mux5~6_combout ),
	.cin(gnd),
	.combout(Mux5),
	.cout());
// synopsys translate_off
defparam \Mux5~9 .lut_mask = 16'hF388;
defparam \Mux5~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N6
cycloneive_lcell_comb \Mux5~19 (
// Equation(s):
// Mux510 = (instruction_D[23] & ((\Mux5~16_combout  & ((\Mux5~18_combout ))) # (!\Mux5~16_combout  & (\Mux5~11_combout )))) # (!instruction_D[23] & (((\Mux5~16_combout ))))

	.dataa(\Mux5~11_combout ),
	.datab(instruction_D_23),
	.datac(\Mux5~18_combout ),
	.datad(\Mux5~16_combout ),
	.cin(gnd),
	.combout(Mux510),
	.cout());
// synopsys translate_off
defparam \Mux5~19 .lut_mask = 16'hF388;
defparam \Mux5~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N8
cycloneive_lcell_comb \Mux6~9 (
// Equation(s):
// Mux6 = (instruction_D[21] & ((\Mux6~6_combout  & (\Mux6~8_combout )) # (!\Mux6~6_combout  & ((\Mux6~1_combout ))))) # (!instruction_D[21] & (((\Mux6~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux6~8_combout ),
	.datac(\Mux6~1_combout ),
	.datad(\Mux6~6_combout ),
	.cin(gnd),
	.combout(Mux6),
	.cout());
// synopsys translate_off
defparam \Mux6~9 .lut_mask = 16'hDDA0;
defparam \Mux6~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N24
cycloneive_lcell_comb \Mux6~19 (
// Equation(s):
// Mux64 = (instruction_D[24] & ((\Mux6~16_combout  & ((\Mux6~18_combout ))) # (!\Mux6~16_combout  & (\Mux6~11_combout )))) # (!instruction_D[24] & (((\Mux6~16_combout ))))

	.dataa(\Mux6~11_combout ),
	.datab(instruction_D_24),
	.datac(\Mux6~16_combout ),
	.datad(\Mux6~18_combout ),
	.cin(gnd),
	.combout(Mux64),
	.cout());
// synopsys translate_off
defparam \Mux6~19 .lut_mask = 16'hF838;
defparam \Mux6~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N18
cycloneive_lcell_comb \Mux7~9 (
// Equation(s):
// Mux7 = (instruction_D[21] & ((\Mux7~6_combout  & (\Mux7~8_combout )) # (!\Mux7~6_combout  & ((\Mux7~1_combout ))))) # (!instruction_D[21] & (((\Mux7~6_combout ))))

	.dataa(\Mux7~8_combout ),
	.datab(instruction_D_21),
	.datac(\Mux7~1_combout ),
	.datad(\Mux7~6_combout ),
	.cin(gnd),
	.combout(Mux7),
	.cout());
// synopsys translate_off
defparam \Mux7~9 .lut_mask = 16'hBBC0;
defparam \Mux7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N8
cycloneive_lcell_comb \Mux7~19 (
// Equation(s):
// Mux71 = (instruction_D[23] & ((\Mux7~16_combout  & ((\Mux7~18_combout ))) # (!\Mux7~16_combout  & (\Mux7~11_combout )))) # (!instruction_D[23] & (((\Mux7~16_combout ))))

	.dataa(\Mux7~11_combout ),
	.datab(instruction_D_23),
	.datac(\Mux7~16_combout ),
	.datad(\Mux7~18_combout ),
	.cin(gnd),
	.combout(Mux71),
	.cout());
// synopsys translate_off
defparam \Mux7~19 .lut_mask = 16'hF838;
defparam \Mux7~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N26
cycloneive_lcell_comb \Mux8~9 (
// Equation(s):
// Mux8 = (instruction_D[21] & ((\Mux8~6_combout  & ((\Mux8~8_combout ))) # (!\Mux8~6_combout  & (\Mux8~1_combout )))) # (!instruction_D[21] & (((\Mux8~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux8~1_combout ),
	.datac(\Mux8~8_combout ),
	.datad(\Mux8~6_combout ),
	.cin(gnd),
	.combout(Mux8),
	.cout());
// synopsys translate_off
defparam \Mux8~9 .lut_mask = 16'hF588;
defparam \Mux8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N30
cycloneive_lcell_comb \Mux8~19 (
// Equation(s):
// Mux81 = (instruction_D[24] & ((\Mux8~16_combout  & (\Mux8~18_combout )) # (!\Mux8~16_combout  & ((\Mux8~11_combout ))))) # (!instruction_D[24] & (((\Mux8~16_combout ))))

	.dataa(instruction_D_24),
	.datab(\Mux8~18_combout ),
	.datac(\Mux8~16_combout ),
	.datad(\Mux8~11_combout ),
	.cin(gnd),
	.combout(Mux81),
	.cout());
// synopsys translate_off
defparam \Mux8~19 .lut_mask = 16'hDAD0;
defparam \Mux8~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N22
cycloneive_lcell_comb \Mux9~9 (
// Equation(s):
// Mux9 = (instruction_D[21] & ((\Mux9~6_combout  & ((\Mux9~8_combout ))) # (!\Mux9~6_combout  & (\Mux9~1_combout )))) # (!instruction_D[21] & (((\Mux9~6_combout ))))

	.dataa(\Mux9~1_combout ),
	.datab(instruction_D_21),
	.datac(\Mux9~8_combout ),
	.datad(\Mux9~6_combout ),
	.cin(gnd),
	.combout(Mux9),
	.cout());
// synopsys translate_off
defparam \Mux9~9 .lut_mask = 16'hF388;
defparam \Mux9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N24
cycloneive_lcell_comb \Mux9~19 (
// Equation(s):
// Mux91 = (instruction_D[23] & ((\Mux9~16_combout  & (\Mux9~18_combout )) # (!\Mux9~16_combout  & ((\Mux9~11_combout ))))) # (!instruction_D[23] & (((\Mux9~16_combout ))))

	.dataa(instruction_D_23),
	.datab(\Mux9~18_combout ),
	.datac(\Mux9~11_combout ),
	.datad(\Mux9~16_combout ),
	.cin(gnd),
	.combout(Mux91),
	.cout());
// synopsys translate_off
defparam \Mux9~19 .lut_mask = 16'hDDA0;
defparam \Mux9~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N2
cycloneive_lcell_comb \Mux10~9 (
// Equation(s):
// Mux10 = (instruction_D[21] & ((\Mux10~6_combout  & ((\Mux10~8_combout ))) # (!\Mux10~6_combout  & (\Mux10~1_combout )))) # (!instruction_D[21] & (((\Mux10~6_combout ))))

	.dataa(\Mux10~1_combout ),
	.datab(instruction_D_21),
	.datac(\Mux10~8_combout ),
	.datad(\Mux10~6_combout ),
	.cin(gnd),
	.combout(Mux10),
	.cout());
// synopsys translate_off
defparam \Mux10~9 .lut_mask = 16'hF388;
defparam \Mux10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N22
cycloneive_lcell_comb \Mux10~19 (
// Equation(s):
// Mux101 = (\Mux10~16_combout  & ((\Mux10~18_combout ) # ((!instruction_D[24])))) # (!\Mux10~16_combout  & (((instruction_D[24] & \Mux10~11_combout ))))

	.dataa(\Mux10~16_combout ),
	.datab(\Mux10~18_combout ),
	.datac(instruction_D_24),
	.datad(\Mux10~11_combout ),
	.cin(gnd),
	.combout(Mux101),
	.cout());
// synopsys translate_off
defparam \Mux10~19 .lut_mask = 16'hDA8A;
defparam \Mux10~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N4
cycloneive_lcell_comb \Mux11~9 (
// Equation(s):
// Mux111 = (instruction_D[21] & ((\Mux11~6_combout  & (\Mux11~8_combout )) # (!\Mux11~6_combout  & ((\Mux11~1_combout ))))) # (!instruction_D[21] & (((\Mux11~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux11~8_combout ),
	.datac(\Mux11~6_combout ),
	.datad(\Mux11~1_combout ),
	.cin(gnd),
	.combout(Mux111),
	.cout());
// synopsys translate_off
defparam \Mux11~9 .lut_mask = 16'hDAD0;
defparam \Mux11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N30
cycloneive_lcell_comb \Mux11~19 (
// Equation(s):
// Mux112 = (instruction_D[23] & ((\Mux11~16_combout  & (\Mux11~18_combout )) # (!\Mux11~16_combout  & ((\Mux11~11_combout ))))) # (!instruction_D[23] & (\Mux11~16_combout ))

	.dataa(instruction_D_23),
	.datab(\Mux11~16_combout ),
	.datac(\Mux11~18_combout ),
	.datad(\Mux11~11_combout ),
	.cin(gnd),
	.combout(Mux112),
	.cout());
// synopsys translate_off
defparam \Mux11~19 .lut_mask = 16'hE6C4;
defparam \Mux11~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N4
cycloneive_lcell_comb \Mux12~9 (
// Equation(s):
// Mux12 = (instruction_D[21] & ((\Mux12~6_combout  & (\Mux12~8_combout )) # (!\Mux12~6_combout  & ((\Mux12~1_combout ))))) # (!instruction_D[21] & (((\Mux12~6_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux12~8_combout ),
	.datac(\Mux12~1_combout ),
	.datad(\Mux12~6_combout ),
	.cin(gnd),
	.combout(Mux12),
	.cout());
// synopsys translate_off
defparam \Mux12~9 .lut_mask = 16'hDDA0;
defparam \Mux12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N8
cycloneive_lcell_comb \Mux12~19 (
// Equation(s):
// Mux121 = (instruction_D[24] & ((\Mux12~16_combout  & (\Mux12~18_combout )) # (!\Mux12~16_combout  & ((\Mux12~11_combout ))))) # (!instruction_D[24] & (((\Mux12~16_combout ))))

	.dataa(\Mux12~18_combout ),
	.datab(instruction_D_24),
	.datac(\Mux12~11_combout ),
	.datad(\Mux12~16_combout ),
	.cin(gnd),
	.combout(Mux121),
	.cout());
// synopsys translate_off
defparam \Mux12~19 .lut_mask = 16'hBBC0;
defparam \Mux12~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N14
cycloneive_lcell_comb \Mux13~9 (
// Equation(s):
// Mux13 = (instruction_D[21] & ((\Mux13~6_combout  & (\Mux13~8_combout )) # (!\Mux13~6_combout  & ((\Mux13~1_combout ))))) # (!instruction_D[21] & (((\Mux13~6_combout ))))

	.dataa(\Mux13~8_combout ),
	.datab(instruction_D_21),
	.datac(\Mux13~1_combout ),
	.datad(\Mux13~6_combout ),
	.cin(gnd),
	.combout(Mux13),
	.cout());
// synopsys translate_off
defparam \Mux13~9 .lut_mask = 16'hBBC0;
defparam \Mux13~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N10
cycloneive_lcell_comb \Mux13~19 (
// Equation(s):
// Mux131 = (instruction_D[23] & ((\Mux13~16_combout  & ((\Mux13~18_combout ))) # (!\Mux13~16_combout  & (\Mux13~11_combout )))) # (!instruction_D[23] & (((\Mux13~16_combout ))))

	.dataa(instruction_D_23),
	.datab(\Mux13~11_combout ),
	.datac(\Mux13~18_combout ),
	.datad(\Mux13~16_combout ),
	.cin(gnd),
	.combout(Mux131),
	.cout());
// synopsys translate_off
defparam \Mux13~19 .lut_mask = 16'hF588;
defparam \Mux13~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N2
cycloneive_lcell_comb \Mux14~9 (
// Equation(s):
// Mux14 = (instruction_D[21] & ((\Mux14~6_combout  & (\Mux14~8_combout )) # (!\Mux14~6_combout  & ((\Mux14~1_combout ))))) # (!instruction_D[21] & (\Mux14~6_combout ))

	.dataa(instruction_D_21),
	.datab(\Mux14~6_combout ),
	.datac(\Mux14~8_combout ),
	.datad(\Mux14~1_combout ),
	.cin(gnd),
	.combout(Mux14),
	.cout());
// synopsys translate_off
defparam \Mux14~9 .lut_mask = 16'hE6C4;
defparam \Mux14~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N8
cycloneive_lcell_comb \Mux14~19 (
// Equation(s):
// Mux141 = (instruction_D[24] & ((\Mux14~16_combout  & ((\Mux14~18_combout ))) # (!\Mux14~16_combout  & (\Mux14~11_combout )))) # (!instruction_D[24] & (((\Mux14~16_combout ))))

	.dataa(\Mux14~11_combout ),
	.datab(instruction_D_24),
	.datac(\Mux14~16_combout ),
	.datad(\Mux14~18_combout ),
	.cin(gnd),
	.combout(Mux141),
	.cout());
// synopsys translate_off
defparam \Mux14~19 .lut_mask = 16'hF838;
defparam \Mux14~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N14
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// Mux311 = (instruction_D[21] & ((\Mux31~6_combout  & ((\Mux31~8_combout ))) # (!\Mux31~6_combout  & (\Mux31~1_combout )))) # (!instruction_D[21] & (((\Mux31~6_combout ))))

	.dataa(\Mux31~1_combout ),
	.datab(instruction_D_21),
	.datac(\Mux31~8_combout ),
	.datad(\Mux31~6_combout ),
	.cin(gnd),
	.combout(Mux311),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'hF388;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N26
cycloneive_lcell_comb \Mux31~19 (
// Equation(s):
// Mux312 = (instruction_D[23] & ((\Mux31~16_combout  & ((\Mux31~18_combout ))) # (!\Mux31~16_combout  & (\Mux31~11_combout )))) # (!instruction_D[23] & (((\Mux31~16_combout ))))

	.dataa(\Mux31~11_combout ),
	.datab(instruction_D_23),
	.datac(\Mux31~18_combout ),
	.datad(\Mux31~16_combout ),
	.cin(gnd),
	.combout(Mux312),
	.cout());
// synopsys translate_off
defparam \Mux31~19 .lut_mask = 16'hF388;
defparam \Mux31~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N20
cycloneive_lcell_comb \Decoder0~2 (
// Equation(s):
// \Decoder0~2_combout  = (!wsel_WB[3] & (!wsel_WB[1] & (\regWrite_WB~q  & wsel_WB[4])))

	.dataa(wsel_WB_3),
	.datab(wsel_WB_1),
	.datac(regWrite_WB),
	.datad(wsel_WB_4),
	.cin(gnd),
	.combout(\Decoder0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~2 .lut_mask = 16'h1000;
defparam \Decoder0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N28
cycloneive_lcell_comb \Decoder0~4 (
// Equation(s):
// \Decoder0~4_combout  = (!wsel_WB[2] & (wsel_WB[0] & \Decoder0~2_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~4 .lut_mask = 16'h5000;
defparam \Decoder0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y28_N5
dffeas \rfile[17][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][31] .is_wysiwyg = "true";
defparam \rfile[17][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N30
cycloneive_lcell_comb \Decoder0~3 (
// Equation(s):
// \Decoder0~3_combout  = (wsel_WB[2] & (wsel_WB[0] & \Decoder0~2_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~3 .lut_mask = 16'hA000;
defparam \Decoder0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N1
dffeas \rfile[21][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][31] .is_wysiwyg = "true";
defparam \rfile[21][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N4
cycloneive_lcell_comb \Mux32~0 (
// Equation(s):
// \Mux32~0_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[21][31]~q ))) # (!instruction_D[18] & (\rfile[17][31]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[17][31]~q ),
	.datad(\rfile[21][31]~q ),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~0 .lut_mask = 16'hDC98;
defparam \Mux32~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N30
cycloneive_lcell_comb \rfile[25][31]~feeder (
// Equation(s):
// \rfile[25][31]~feeder_combout  = \wdat_WB[31]~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_31),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[25][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[25][31]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[25][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N4
cycloneive_lcell_comb \Decoder0~0 (
// Equation(s):
// \Decoder0~0_combout  = (wsel_WB[4] & (wsel_WB[3] & (!wsel_WB[1] & \regWrite_WB~q )))

	.dataa(wsel_WB_4),
	.datab(wsel_WB_3),
	.datac(wsel_WB_1),
	.datad(regWrite_WB),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~0 .lut_mask = 16'h0800;
defparam \Decoder0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N2
cycloneive_lcell_comb \Decoder0~1 (
// Equation(s):
// \Decoder0~1_combout  = (wsel_WB[0] & (\Decoder0~0_combout  & !wsel_WB[2]))

	.dataa(gnd),
	.datab(wsel_WB_0),
	.datac(\Decoder0~0_combout ),
	.datad(wsel_WB_2),
	.cin(gnd),
	.combout(\Decoder0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~1 .lut_mask = 16'h00C0;
defparam \Decoder0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N31
dffeas \rfile[25][31] (
	.clk(!CLK),
	.d(\rfile[25][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][31] .is_wysiwyg = "true";
defparam \rfile[25][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N20
cycloneive_lcell_comb \Decoder0~5 (
// Equation(s):
// \Decoder0~5_combout  = (wsel_WB[0] & (\Decoder0~0_combout  & wsel_WB[2]))

	.dataa(gnd),
	.datab(wsel_WB_0),
	.datac(\Decoder0~0_combout ),
	.datad(wsel_WB_2),
	.cin(gnd),
	.combout(\Decoder0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~5 .lut_mask = 16'hC000;
defparam \Decoder0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N7
dffeas \rfile[29][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][31] .is_wysiwyg = "true";
defparam \rfile[29][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N8
cycloneive_lcell_comb \Mux32~1 (
// Equation(s):
// \Mux32~1_combout  = (\Mux32~0_combout  & (((\rfile[29][31]~q )) # (!instruction_D[19]))) # (!\Mux32~0_combout  & (instruction_D[19] & (\rfile[25][31]~q )))

	.dataa(\Mux32~0_combout ),
	.datab(instruction_D_19),
	.datac(\rfile[25][31]~q ),
	.datad(\rfile[29][31]~q ),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~1 .lut_mask = 16'hEA62;
defparam \Mux32~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N28
cycloneive_lcell_comb \Decoder0~8 (
// Equation(s):
// \Decoder0~8_combout  = (wsel_WB[4] & (wsel_WB[3] & (wsel_WB[1] & \regWrite_WB~q )))

	.dataa(wsel_WB_4),
	.datab(wsel_WB_3),
	.datac(wsel_WB_1),
	.datad(regWrite_WB),
	.cin(gnd),
	.combout(\Decoder0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~8 .lut_mask = 16'h8000;
defparam \Decoder0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N6
cycloneive_lcell_comb \Decoder0~16 (
// Equation(s):
// \Decoder0~16_combout  = (!wsel_WB[2] & (wsel_WB[0] & \Decoder0~8_combout ))

	.dataa(wsel_WB_2),
	.datab(wsel_WB_0),
	.datac(gnd),
	.datad(\Decoder0~8_combout ),
	.cin(gnd),
	.combout(\Decoder0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~16 .lut_mask = 16'h4400;
defparam \Decoder0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N5
dffeas \rfile[27][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][31] .is_wysiwyg = "true";
defparam \rfile[27][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N18
cycloneive_lcell_comb \Decoder0~6 (
// Equation(s):
// \Decoder0~6_combout  = (wsel_WB[4] & (wsel_WB[1] & (!wsel_WB[3] & \regWrite_WB~q )))

	.dataa(wsel_WB_4),
	.datab(wsel_WB_1),
	.datac(wsel_WB_3),
	.datad(regWrite_WB),
	.cin(gnd),
	.combout(\Decoder0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~6 .lut_mask = 16'h0800;
defparam \Decoder0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N6
cycloneive_lcell_comb \Decoder0~17 (
// Equation(s):
// \Decoder0~17_combout  = (wsel_WB[2] & (wsel_WB[0] & \Decoder0~6_combout ))

	.dataa(gnd),
	.datab(wsel_WB_2),
	.datac(wsel_WB_0),
	.datad(\Decoder0~6_combout ),
	.cin(gnd),
	.combout(\Decoder0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~17 .lut_mask = 16'hC000;
defparam \Decoder0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y31_N21
dffeas \rfile[23][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][31] .is_wysiwyg = "true";
defparam \rfile[23][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N12
cycloneive_lcell_comb \rfile[19][31]~feeder (
// Equation(s):
// \rfile[19][31]~feeder_combout  = \wdat_WB[31]~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_31),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[19][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[19][31]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[19][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N20
cycloneive_lcell_comb \Decoder0~18 (
// Equation(s):
// \Decoder0~18_combout  = (!wsel_WB[2] & (wsel_WB[0] & \Decoder0~6_combout ))

	.dataa(gnd),
	.datab(wsel_WB_2),
	.datac(wsel_WB_0),
	.datad(\Decoder0~6_combout ),
	.cin(gnd),
	.combout(\Decoder0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~18 .lut_mask = 16'h3000;
defparam \Decoder0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y28_N13
dffeas \rfile[19][31] (
	.clk(!CLK),
	.d(\rfile[19][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][31] .is_wysiwyg = "true";
defparam \rfile[19][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N20
cycloneive_lcell_comb \Mux32~7 (
// Equation(s):
// \Mux32~7_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[23][31]~q )) # (!instruction_D[18] & ((\rfile[19][31]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[23][31]~q ),
	.datad(\rfile[19][31]~q ),
	.cin(gnd),
	.combout(\Mux32~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~7 .lut_mask = 16'hD9C8;
defparam \Mux32~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N22
cycloneive_lcell_comb \rfile[31][31]~feeder (
// Equation(s):
// \rfile[31][31]~feeder_combout  = \wdat_WB[31]~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_31),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[31][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[31][31]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[31][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N26
cycloneive_lcell_comb \Decoder0~19 (
// Equation(s):
// \Decoder0~19_combout  = (wsel_WB[2] & (wsel_WB[0] & \Decoder0~8_combout ))

	.dataa(wsel_WB_2),
	.datab(wsel_WB_0),
	.datac(gnd),
	.datad(\Decoder0~8_combout ),
	.cin(gnd),
	.combout(\Decoder0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~19 .lut_mask = 16'h8800;
defparam \Decoder0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N23
dffeas \rfile[31][31] (
	.clk(!CLK),
	.d(\rfile[31][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][31] .is_wysiwyg = "true";
defparam \rfile[31][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N12
cycloneive_lcell_comb \Mux32~8 (
// Equation(s):
// \Mux32~8_combout  = (instruction_D[19] & ((\Mux32~7_combout  & ((\rfile[31][31]~q ))) # (!\Mux32~7_combout  & (\rfile[27][31]~q )))) # (!instruction_D[19] & (((\Mux32~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[27][31]~q ),
	.datac(\Mux32~7_combout ),
	.datad(\rfile[31][31]~q ),
	.cin(gnd),
	.combout(\Mux32~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~8 .lut_mask = 16'hF858;
defparam \Mux32~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N0
cycloneive_lcell_comb \rfile[28][31]~feeder (
// Equation(s):
// \rfile[28][31]~feeder_combout  = \wdat_WB[31]~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_31),
	.cin(gnd),
	.combout(\rfile[28][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][31]~feeder .lut_mask = 16'hFF00;
defparam \rfile[28][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N16
cycloneive_lcell_comb \Decoder0~15 (
// Equation(s):
// \Decoder0~15_combout  = (wsel_WB[2] & (!wsel_WB[0] & \Decoder0~0_combout ))

	.dataa(gnd),
	.datab(wsel_WB_2),
	.datac(wsel_WB_0),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~15 .lut_mask = 16'h0C00;
defparam \Decoder0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y32_N1
dffeas \rfile[28][31] (
	.clk(!CLK),
	.d(\rfile[28][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][31] .is_wysiwyg = "true";
defparam \rfile[28][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N14
cycloneive_lcell_comb \Decoder0~13 (
// Equation(s):
// \Decoder0~13_combout  = (!wsel_WB[2] & (!wsel_WB[0] & \Decoder0~0_combout ))

	.dataa(gnd),
	.datab(wsel_WB_2),
	.datac(wsel_WB_0),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~13 .lut_mask = 16'h0300;
defparam \Decoder0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y33_N9
dffeas \rfile[24][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][31] .is_wysiwyg = "true";
defparam \rfile[24][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N14
cycloneive_lcell_comb \Decoder0~14 (
// Equation(s):
// \Decoder0~14_combout  = (!wsel_WB[0] & (\Decoder0~2_combout  & !wsel_WB[2]))

	.dataa(gnd),
	.datab(wsel_WB_0),
	.datac(\Decoder0~2_combout ),
	.datad(wsel_WB_2),
	.cin(gnd),
	.combout(\Decoder0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~14 .lut_mask = 16'h0030;
defparam \Decoder0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y33_N19
dffeas \rfile[16][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][31] .is_wysiwyg = "true";
defparam \rfile[16][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N18
cycloneive_lcell_comb \Mux32~4 (
// Equation(s):
// \Mux32~4_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[24][31]~q )) # (!instruction_D[19] & ((\rfile[16][31]~q )))))

	.dataa(instruction_D_18),
	.datab(\rfile[24][31]~q ),
	.datac(\rfile[16][31]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~4 .lut_mask = 16'hEE50;
defparam \Mux32~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N18
cycloneive_lcell_comb \Mux32~5 (
// Equation(s):
// \Mux32~5_combout  = (instruction_D[18] & ((\Mux32~4_combout  & ((\rfile[28][31]~q ))) # (!\Mux32~4_combout  & (\rfile[20][31]~q )))) # (!instruction_D[18] & (((\Mux32~4_combout ))))

	.dataa(\rfile[20][31]~q ),
	.datab(\rfile[28][31]~q ),
	.datac(instruction_D_18),
	.datad(\Mux32~4_combout ),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~5 .lut_mask = 16'hCFA0;
defparam \Mux32~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N26
cycloneive_lcell_comb \Decoder0~7 (
// Equation(s):
// \Decoder0~7_combout  = (wsel_WB[2] & (!wsel_WB[0] & \Decoder0~6_combout ))

	.dataa(wsel_WB_2),
	.datab(wsel_WB_0),
	.datac(gnd),
	.datad(\Decoder0~6_combout ),
	.cin(gnd),
	.combout(\Decoder0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~7 .lut_mask = 16'h2200;
defparam \Decoder0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y34_N5
dffeas \rfile[22][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][31] .is_wysiwyg = "true";
defparam \rfile[22][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N4
cycloneive_lcell_comb \Decoder0~11 (
// Equation(s):
// \Decoder0~11_combout  = (!wsel_WB[0] & (wsel_WB[2] & \Decoder0~8_combout ))

	.dataa(wsel_WB_0),
	.datab(wsel_WB_2),
	.datac(gnd),
	.datad(\Decoder0~8_combout ),
	.cin(gnd),
	.combout(\Decoder0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~11 .lut_mask = 16'h4400;
defparam \Decoder0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y36_N15
dffeas \rfile[30][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][31] .is_wysiwyg = "true";
defparam \rfile[30][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N4
cycloneive_lcell_comb \Mux32~3 (
// Equation(s):
// \Mux32~3_combout  = (\Mux32~2_combout  & (((\rfile[30][31]~q )) # (!instruction_D[18]))) # (!\Mux32~2_combout  & (instruction_D[18] & (\rfile[22][31]~q )))

	.dataa(\Mux32~2_combout ),
	.datab(instruction_D_18),
	.datac(\rfile[22][31]~q ),
	.datad(\rfile[30][31]~q ),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~3 .lut_mask = 16'hEA62;
defparam \Mux32~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N10
cycloneive_lcell_comb \Mux32~6 (
// Equation(s):
// \Mux32~6_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & ((\Mux32~3_combout ))) # (!instruction_D[17] & (\Mux32~5_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux32~5_combout ),
	.datac(instruction_D_17),
	.datad(\Mux32~3_combout ),
	.cin(gnd),
	.combout(\Mux32~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~6 .lut_mask = 16'hF4A4;
defparam \Mux32~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N8
cycloneive_lcell_comb \rfile[11][31]~feeder (
// Equation(s):
// \rfile[11][31]~feeder_combout  = \wdat_WB[31]~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_31),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[11][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][31]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[11][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N24
cycloneive_lcell_comb \Decoder0~22 (
// Equation(s):
// \Decoder0~22_combout  = (\regWrite_WB~q  & (wsel_WB[3] & (!wsel_WB[4] & wsel_WB[1])))

	.dataa(regWrite_WB),
	.datab(wsel_WB_3),
	.datac(wsel_WB_4),
	.datad(wsel_WB_1),
	.cin(gnd),
	.combout(\Decoder0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~22 .lut_mask = 16'h0800;
defparam \Decoder0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N24
cycloneive_lcell_comb \Decoder0~25 (
// Equation(s):
// \Decoder0~25_combout  = (!wsel_WB[2] & (wsel_WB[0] & \Decoder0~22_combout ))

	.dataa(wsel_WB_2),
	.datab(wsel_WB_0),
	.datac(gnd),
	.datad(\Decoder0~22_combout ),
	.cin(gnd),
	.combout(\Decoder0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~25 .lut_mask = 16'h4400;
defparam \Decoder0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N9
dffeas \rfile[11][31] (
	.clk(!CLK),
	.d(\rfile[11][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][31] .is_wysiwyg = "true";
defparam \rfile[11][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N10
cycloneive_lcell_comb \Decoder0~23 (
// Equation(s):
// \Decoder0~23_combout  = (!wsel_WB[2] & (!wsel_WB[0] & \Decoder0~22_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~22_combout ),
	.cin(gnd),
	.combout(\Decoder0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~23 .lut_mask = 16'h0500;
defparam \Decoder0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N29
dffeas \rfile[10][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][31] .is_wysiwyg = "true";
defparam \rfile[10][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N28
cycloneive_lcell_comb \Mux32~10 (
// Equation(s):
// \Mux32~10_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][31]~q ))) # (!instruction_D[17] & (\rfile[8][31]~q ))))

	.dataa(\rfile[8][31]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[10][31]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux32~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~10 .lut_mask = 16'hFC22;
defparam \Mux32~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N24
cycloneive_lcell_comb \rfile[9][31]~feeder (
// Equation(s):
// \rfile[9][31]~feeder_combout  = \wdat_WB[31]~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_31),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[9][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][31]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[9][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N2
cycloneive_lcell_comb \Decoder0~20 (
// Equation(s):
// \Decoder0~20_combout  = (!wsel_WB[4] & (!wsel_WB[1] & (wsel_WB[3] & \regWrite_WB~q )))

	.dataa(wsel_WB_4),
	.datab(wsel_WB_1),
	.datac(wsel_WB_3),
	.datad(regWrite_WB),
	.cin(gnd),
	.combout(\Decoder0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~20 .lut_mask = 16'h1000;
defparam \Decoder0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N24
cycloneive_lcell_comb \Decoder0~21 (
// Equation(s):
// \Decoder0~21_combout  = (wsel_WB[0] & (\Decoder0~20_combout  & !wsel_WB[2]))

	.dataa(wsel_WB_0),
	.datab(\Decoder0~20_combout ),
	.datac(wsel_WB_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~21 .lut_mask = 16'h0808;
defparam \Decoder0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N25
dffeas \rfile[9][31] (
	.clk(!CLK),
	.d(\rfile[9][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][31] .is_wysiwyg = "true";
defparam \rfile[9][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N20
cycloneive_lcell_comb \Mux32~11 (
// Equation(s):
// \Mux32~11_combout  = (instruction_D[16] & ((\Mux32~10_combout  & (\rfile[11][31]~q )) # (!\Mux32~10_combout  & ((\rfile[9][31]~q ))))) # (!instruction_D[16] & (((\Mux32~10_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][31]~q ),
	.datac(\Mux32~10_combout ),
	.datad(\rfile[9][31]~q ),
	.cin(gnd),
	.combout(\Mux32~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~11 .lut_mask = 16'hDAD0;
defparam \Mux32~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N16
cycloneive_lcell_comb \Decoder0~26 (
// Equation(s):
// \Decoder0~26_combout  = (\regWrite_WB~q  & (!wsel_WB[3] & (!wsel_WB[4] & wsel_WB[1])))

	.dataa(regWrite_WB),
	.datab(wsel_WB_3),
	.datac(wsel_WB_4),
	.datad(wsel_WB_1),
	.cin(gnd),
	.combout(\Decoder0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~26 .lut_mask = 16'h0200;
defparam \Decoder0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N14
cycloneive_lcell_comb \Decoder0~27 (
// Equation(s):
// \Decoder0~27_combout  = (wsel_WB[2] & (!wsel_WB[0] & \Decoder0~26_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~26_combout ),
	.cin(gnd),
	.combout(\Decoder0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~27 .lut_mask = 16'h0A00;
defparam \Decoder0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N17
dffeas \rfile[6][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][31] .is_wysiwyg = "true";
defparam \rfile[6][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N28
cycloneive_lcell_comb \Decoder0~28 (
// Equation(s):
// \Decoder0~28_combout  = (\regWrite_WB~q  & (!wsel_WB[3] & (!wsel_WB[4] & !wsel_WB[1])))

	.dataa(regWrite_WB),
	.datab(wsel_WB_3),
	.datac(wsel_WB_4),
	.datad(wsel_WB_1),
	.cin(gnd),
	.combout(\Decoder0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~28 .lut_mask = 16'h0002;
defparam \Decoder0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N6
cycloneive_lcell_comb \Decoder0~29 (
// Equation(s):
// \Decoder0~29_combout  = (wsel_WB[2] & (wsel_WB[0] & \Decoder0~28_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~28_combout ),
	.cin(gnd),
	.combout(\Decoder0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~29 .lut_mask = 16'hA000;
defparam \Decoder0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N13
dffeas \rfile[5][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][31] .is_wysiwyg = "true";
defparam \rfile[5][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N12
cycloneive_lcell_comb \Mux32~12 (
// Equation(s):
// \Mux32~12_combout  = (instruction_D[17] & (((instruction_D[16])))) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][31]~q ))) # (!instruction_D[16] & (\rfile[4][31]~q ))))

	.dataa(\rfile[4][31]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[5][31]~q ),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux32~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~12 .lut_mask = 16'hFC22;
defparam \Mux32~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N16
cycloneive_lcell_comb \Mux32~13 (
// Equation(s):
// \Mux32~13_combout  = (instruction_D[17] & ((\Mux32~12_combout  & (\rfile[7][31]~q )) # (!\Mux32~12_combout  & ((\rfile[6][31]~q ))))) # (!instruction_D[17] & (((\Mux32~12_combout ))))

	.dataa(\rfile[7][31]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[6][31]~q ),
	.datad(\Mux32~12_combout ),
	.cin(gnd),
	.combout(\Mux32~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~13 .lut_mask = 16'hBBC0;
defparam \Mux32~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N26
cycloneive_lcell_comb \Decoder0~34 (
// Equation(s):
// \Decoder0~34_combout  = (!wsel_WB[2] & (!wsel_WB[0] & \Decoder0~26_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~26_combout ),
	.cin(gnd),
	.combout(\Decoder0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~34 .lut_mask = 16'h0500;
defparam \Decoder0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N19
dffeas \rfile[2][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][31] .is_wysiwyg = "true";
defparam \rfile[2][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N8
cycloneive_lcell_comb \Decoder0~32 (
// Equation(s):
// \Decoder0~32_combout  = (wsel_WB[0] & (!wsel_WB[2] & \Decoder0~26_combout ))

	.dataa(wsel_WB_0),
	.datab(wsel_WB_2),
	.datac(gnd),
	.datad(\Decoder0~26_combout ),
	.cin(gnd),
	.combout(\Decoder0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~32 .lut_mask = 16'h2200;
defparam \Decoder0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y34_N17
dffeas \rfile[3][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][31] .is_wysiwyg = "true";
defparam \rfile[3][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N0
cycloneive_lcell_comb \Decoder0~33 (
// Equation(s):
// \Decoder0~33_combout  = (!wsel_WB[2] & (wsel_WB[0] & \Decoder0~28_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~28_combout ),
	.cin(gnd),
	.combout(\Decoder0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~33 .lut_mask = 16'h5000;
defparam \Decoder0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y34_N15
dffeas \rfile[1][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][31] .is_wysiwyg = "true";
defparam \rfile[1][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N16
cycloneive_lcell_comb \Mux32~14 (
// Equation(s):
// \Mux32~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][31]~q )) # (!instruction_D[17] & ((\rfile[1][31]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[3][31]~q ),
	.datad(\rfile[1][31]~q ),
	.cin(gnd),
	.combout(\Mux32~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~14 .lut_mask = 16'hA280;
defparam \Mux32~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N18
cycloneive_lcell_comb \Mux32~15 (
// Equation(s):
// \Mux32~15_combout  = (\Mux32~14_combout ) # ((!instruction_D[16] & (instruction_D[17] & \rfile[2][31]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[2][31]~q ),
	.datad(\Mux32~14_combout ),
	.cin(gnd),
	.combout(\Mux32~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~15 .lut_mask = 16'hFF40;
defparam \Mux32~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N8
cycloneive_lcell_comb \Mux32~16 (
// Equation(s):
// \Mux32~16_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\Mux32~13_combout )) # (!instruction_D[18] & ((\Mux32~15_combout )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux32~13_combout ),
	.datad(\Mux32~15_combout ),
	.cin(gnd),
	.combout(\Mux32~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~16 .lut_mask = 16'hD9C8;
defparam \Mux32~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N12
cycloneive_lcell_comb \rfile[14][31]~feeder (
// Equation(s):
// \rfile[14][31]~feeder_combout  = \wdat_WB[31]~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_31),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[14][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][31]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[14][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N26
cycloneive_lcell_comb \Decoder0~35 (
// Equation(s):
// \Decoder0~35_combout  = (wsel_WB[2] & (!wsel_WB[0] & \Decoder0~22_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~22_combout ),
	.cin(gnd),
	.combout(\Decoder0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~35 .lut_mask = 16'h0A00;
defparam \Decoder0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N13
dffeas \rfile[14][31] (
	.clk(!CLK),
	.d(\rfile[14][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][31] .is_wysiwyg = "true";
defparam \rfile[14][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N18
cycloneive_lcell_comb \Decoder0~38 (
// Equation(s):
// \Decoder0~38_combout  = (wsel_WB[2] & (wsel_WB[0] & \Decoder0~22_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~22_combout ),
	.cin(gnd),
	.combout(\Decoder0~38_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~38 .lut_mask = 16'hA000;
defparam \Decoder0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N27
dffeas \rfile[15][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][31] .is_wysiwyg = "true";
defparam \rfile[15][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N22
cycloneive_lcell_comb \Decoder0~37 (
// Equation(s):
// \Decoder0~37_combout  = (!wsel_WB[0] & (wsel_WB[2] & \Decoder0~20_combout ))

	.dataa(wsel_WB_0),
	.datab(wsel_WB_2),
	.datac(gnd),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~37_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~37 .lut_mask = 16'h4400;
defparam \Decoder0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N29
dffeas \rfile[12][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][31] .is_wysiwyg = "true";
defparam \rfile[12][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N12
cycloneive_lcell_comb \Decoder0~36 (
// Equation(s):
// \Decoder0~36_combout  = (wsel_WB[2] & (wsel_WB[0] & \Decoder0~20_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~36 .lut_mask = 16'hA000;
defparam \Decoder0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N5
dffeas \rfile[13][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][31] .is_wysiwyg = "true";
defparam \rfile[13][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N28
cycloneive_lcell_comb \Mux32~17 (
// Equation(s):
// \Mux32~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][31]~q ))) # (!instruction_D[16] & (\rfile[12][31]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][31]~q ),
	.datad(\rfile[13][31]~q ),
	.cin(gnd),
	.combout(\Mux32~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~17 .lut_mask = 16'hDC98;
defparam \Mux32~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N26
cycloneive_lcell_comb \Mux32~18 (
// Equation(s):
// \Mux32~18_combout  = (instruction_D[17] & ((\Mux32~17_combout  & ((\rfile[15][31]~q ))) # (!\Mux32~17_combout  & (\rfile[14][31]~q )))) # (!instruction_D[17] & (((\Mux32~17_combout ))))

	.dataa(\rfile[14][31]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[15][31]~q ),
	.datad(\Mux32~17_combout ),
	.cin(gnd),
	.combout(\Mux32~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~18 .lut_mask = 16'hF388;
defparam \Mux32~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N17
dffeas \rfile[21][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][30] .is_wysiwyg = "true";
defparam \rfile[21][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N3
dffeas \rfile[29][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][30] .is_wysiwyg = "true";
defparam \rfile[29][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N9
dffeas \rfile[25][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][30] .is_wysiwyg = "true";
defparam \rfile[25][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N19
dffeas \rfile[17][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][30] .is_wysiwyg = "true";
defparam \rfile[17][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N8
cycloneive_lcell_comb \Mux33~0 (
// Equation(s):
// \Mux33~0_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[25][30]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[17][30]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[25][30]~q ),
	.datad(\rfile[17][30]~q ),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~0 .lut_mask = 16'hB9A8;
defparam \Mux33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N2
cycloneive_lcell_comb \Mux33~1 (
// Equation(s):
// \Mux33~1_combout  = (instruction_D[18] & ((\Mux33~0_combout  & ((\rfile[29][30]~q ))) # (!\Mux33~0_combout  & (\rfile[21][30]~q )))) # (!instruction_D[18] & (((\Mux33~0_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[21][30]~q ),
	.datac(\rfile[29][30]~q ),
	.datad(\Mux33~0_combout ),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~1 .lut_mask = 16'hF588;
defparam \Mux33~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N31
dffeas \rfile[31][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][30] .is_wysiwyg = "true";
defparam \rfile[31][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N5
dffeas \rfile[23][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][30] .is_wysiwyg = "true";
defparam \rfile[23][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N15
dffeas \rfile[19][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][30] .is_wysiwyg = "true";
defparam \rfile[19][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N21
dffeas \rfile[27][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][30] .is_wysiwyg = "true";
defparam \rfile[27][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N20
cycloneive_lcell_comb \Mux33~7 (
// Equation(s):
// \Mux33~7_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[27][30]~q ))) # (!instruction_D[19] & (\rfile[19][30]~q ))))

	.dataa(instruction_D_18),
	.datab(\rfile[19][30]~q ),
	.datac(\rfile[27][30]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux33~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~7 .lut_mask = 16'hFA44;
defparam \Mux33~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N4
cycloneive_lcell_comb \Mux33~8 (
// Equation(s):
// \Mux33~8_combout  = (instruction_D[18] & ((\Mux33~7_combout  & (\rfile[31][30]~q )) # (!\Mux33~7_combout  & ((\rfile[23][30]~q ))))) # (!instruction_D[18] & (((\Mux33~7_combout ))))

	.dataa(\rfile[31][30]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[23][30]~q ),
	.datad(\Mux33~7_combout ),
	.cin(gnd),
	.combout(\Mux33~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~8 .lut_mask = 16'hBBC0;
defparam \Mux33~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N6
cycloneive_lcell_comb \Decoder0~9 (
// Equation(s):
// \Decoder0~9_combout  = (!wsel_WB[0] & (!wsel_WB[2] & \Decoder0~8_combout ))

	.dataa(wsel_WB_0),
	.datab(gnd),
	.datac(wsel_WB_2),
	.datad(\Decoder0~8_combout ),
	.cin(gnd),
	.combout(\Decoder0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~9 .lut_mask = 16'h0500;
defparam \Decoder0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y34_N29
dffeas \rfile[26][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][30] .is_wysiwyg = "true";
defparam \rfile[26][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y34_N11
dffeas \rfile[30][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][30] .is_wysiwyg = "true";
defparam \rfile[30][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N28
cycloneive_lcell_comb \Mux33~3 (
// Equation(s):
// \Mux33~3_combout  = (\Mux33~2_combout  & (((\rfile[30][30]~q )) # (!instruction_D[19]))) # (!\Mux33~2_combout  & (instruction_D[19] & (\rfile[26][30]~q )))

	.dataa(\Mux33~2_combout ),
	.datab(instruction_D_19),
	.datac(\rfile[26][30]~q ),
	.datad(\rfile[30][30]~q ),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~3 .lut_mask = 16'hEA62;
defparam \Mux33~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N9
dffeas \rfile[24][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][30] .is_wysiwyg = "true";
defparam \rfile[24][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N20
cycloneive_lcell_comb \Decoder0~12 (
// Equation(s):
// \Decoder0~12_combout  = (!wsel_WB[0] & (\Decoder0~2_combout  & wsel_WB[2]))

	.dataa(gnd),
	.datab(wsel_WB_0),
	.datac(\Decoder0~2_combout ),
	.datad(wsel_WB_2),
	.cin(gnd),
	.combout(\Decoder0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~12 .lut_mask = 16'h3000;
defparam \Decoder0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y31_N17
dffeas \rfile[20][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][30] .is_wysiwyg = "true";
defparam \rfile[20][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y31_N11
dffeas \rfile[16][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][30] .is_wysiwyg = "true";
defparam \rfile[16][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N16
cycloneive_lcell_comb \Mux33~4 (
// Equation(s):
// \Mux33~4_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[20][30]~q )))) # (!instruction_D[18] & (!instruction_D[19] & ((\rfile[16][30]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[20][30]~q ),
	.datad(\rfile[16][30]~q ),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~4 .lut_mask = 16'hB9A8;
defparam \Mux33~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N8
cycloneive_lcell_comb \Mux33~5 (
// Equation(s):
// \Mux33~5_combout  = (instruction_D[19] & ((\Mux33~4_combout  & (\rfile[28][30]~q )) # (!\Mux33~4_combout  & ((\rfile[24][30]~q ))))) # (!instruction_D[19] & (((\Mux33~4_combout ))))

	.dataa(\rfile[28][30]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[24][30]~q ),
	.datad(\Mux33~4_combout ),
	.cin(gnd),
	.combout(\Mux33~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~5 .lut_mask = 16'hBBC0;
defparam \Mux33~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N20
cycloneive_lcell_comb \Mux33~6 (
// Equation(s):
// \Mux33~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\Mux33~3_combout )) # (!instruction_D[17] & ((\Mux33~5_combout )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux33~3_combout ),
	.datad(\Mux33~5_combout ),
	.cin(gnd),
	.combout(\Mux33~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~6 .lut_mask = 16'hD9C8;
defparam \Mux33~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N1
dffeas \rfile[14][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][30] .is_wysiwyg = "true";
defparam \rfile[14][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N31
dffeas \rfile[15][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][30] .is_wysiwyg = "true";
defparam \rfile[15][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N23
dffeas \rfile[13][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][30] .is_wysiwyg = "true";
defparam \rfile[13][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N25
dffeas \rfile[12][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][30] .is_wysiwyg = "true";
defparam \rfile[12][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N22
cycloneive_lcell_comb \Mux33~17 (
// Equation(s):
// \Mux33~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][30]~q )))) # (!instruction_D[16] & (!instruction_D[17] & ((\rfile[12][30]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[13][30]~q ),
	.datad(\rfile[12][30]~q ),
	.cin(gnd),
	.combout(\Mux33~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~17 .lut_mask = 16'hB9A8;
defparam \Mux33~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N30
cycloneive_lcell_comb \Mux33~18 (
// Equation(s):
// \Mux33~18_combout  = (instruction_D[17] & ((\Mux33~17_combout  & ((\rfile[15][30]~q ))) # (!\Mux33~17_combout  & (\rfile[14][30]~q )))) # (!instruction_D[17] & (((\Mux33~17_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[14][30]~q ),
	.datac(\rfile[15][30]~q ),
	.datad(\Mux33~17_combout ),
	.cin(gnd),
	.combout(\Mux33~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~18 .lut_mask = 16'hF588;
defparam \Mux33~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N28
cycloneive_lcell_comb \rfile[2][30]~feeder (
// Equation(s):
// \rfile[2][30]~feeder_combout  = \wdat_WB[30]~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_30),
	.cin(gnd),
	.combout(\rfile[2][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][30]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N29
dffeas \rfile[2][30] (
	.clk(!CLK),
	.d(\rfile[2][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][30] .is_wysiwyg = "true";
defparam \rfile[2][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y34_N25
dffeas \rfile[3][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][30] .is_wysiwyg = "true";
defparam \rfile[3][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y34_N7
dffeas \rfile[1][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][30] .is_wysiwyg = "true";
defparam \rfile[1][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N24
cycloneive_lcell_comb \Mux33~14 (
// Equation(s):
// \Mux33~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][30]~q )) # (!instruction_D[17] & ((\rfile[1][30]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[3][30]~q ),
	.datad(\rfile[1][30]~q ),
	.cin(gnd),
	.combout(\Mux33~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~14 .lut_mask = 16'hA280;
defparam \Mux33~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N30
cycloneive_lcell_comb \Mux33~15 (
// Equation(s):
// \Mux33~15_combout  = (\Mux33~14_combout ) # ((!instruction_D[16] & (\rfile[2][30]~q  & instruction_D[17])))

	.dataa(instruction_D_16),
	.datab(\rfile[2][30]~q ),
	.datac(instruction_D_17),
	.datad(\Mux33~14_combout ),
	.cin(gnd),
	.combout(\Mux33~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~15 .lut_mask = 16'hFF40;
defparam \Mux33~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N9
dffeas \rfile[9][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][30] .is_wysiwyg = "true";
defparam \rfile[9][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N26
cycloneive_lcell_comb \Decoder0~24 (
// Equation(s):
// \Decoder0~24_combout  = (!wsel_WB[2] & (!wsel_WB[0] & \Decoder0~20_combout ))

	.dataa(gnd),
	.datab(wsel_WB_2),
	.datac(wsel_WB_0),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~24 .lut_mask = 16'h0300;
defparam \Decoder0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N3
dffeas \rfile[8][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][30] .is_wysiwyg = "true";
defparam \rfile[8][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N25
dffeas \rfile[10][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][30] .is_wysiwyg = "true";
defparam \rfile[10][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N2
cycloneive_lcell_comb \Mux33~12 (
// Equation(s):
// \Mux33~12_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][30]~q )))) # (!instruction_D[17] & (!instruction_D[16] & (\rfile[8][30]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[8][30]~q ),
	.datad(\rfile[10][30]~q ),
	.cin(gnd),
	.combout(\Mux33~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~12 .lut_mask = 16'hBA98;
defparam \Mux33~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N8
cycloneive_lcell_comb \Mux33~13 (
// Equation(s):
// \Mux33~13_combout  = (instruction_D[16] & ((\Mux33~12_combout  & (\rfile[11][30]~q )) # (!\Mux33~12_combout  & ((\rfile[9][30]~q ))))) # (!instruction_D[16] & (((\Mux33~12_combout ))))

	.dataa(\rfile[11][30]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[9][30]~q ),
	.datad(\Mux33~12_combout ),
	.cin(gnd),
	.combout(\Mux33~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~13 .lut_mask = 16'hBBC0;
defparam \Mux33~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N22
cycloneive_lcell_comb \Mux33~16 (
// Equation(s):
// \Mux33~16_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\Mux33~13_combout )))) # (!instruction_D[19] & (!instruction_D[18] & (\Mux33~15_combout )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux33~15_combout ),
	.datad(\Mux33~13_combout ),
	.cin(gnd),
	.combout(\Mux33~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~16 .lut_mask = 16'hBA98;
defparam \Mux33~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N1
dffeas \rfile[5][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][30] .is_wysiwyg = "true";
defparam \rfile[5][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N0
cycloneive_lcell_comb \Mux33~10 (
// Equation(s):
// \Mux33~10_combout  = (instruction_D[17] & (((instruction_D[16])))) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][30]~q ))) # (!instruction_D[16] & (\rfile[4][30]~q ))))

	.dataa(\rfile[4][30]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[5][30]~q ),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux33~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~10 .lut_mask = 16'hFC22;
defparam \Mux33~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N25
dffeas \rfile[6][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][30] .is_wysiwyg = "true";
defparam \rfile[6][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N2
cycloneive_lcell_comb \Decoder0~31 (
// Equation(s):
// \Decoder0~31_combout  = (wsel_WB[2] & (wsel_WB[0] & \Decoder0~26_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~26_combout ),
	.cin(gnd),
	.combout(\Decoder0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~31 .lut_mask = 16'hA000;
defparam \Decoder0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N3
dffeas \rfile[7][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][30] .is_wysiwyg = "true";
defparam \rfile[7][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N24
cycloneive_lcell_comb \Mux33~11 (
// Equation(s):
// \Mux33~11_combout  = (instruction_D[17] & ((\Mux33~10_combout  & ((\rfile[7][30]~q ))) # (!\Mux33~10_combout  & (\rfile[6][30]~q )))) # (!instruction_D[17] & (\Mux33~10_combout ))

	.dataa(instruction_D_17),
	.datab(\Mux33~10_combout ),
	.datac(\rfile[6][30]~q ),
	.datad(\rfile[7][30]~q ),
	.cin(gnd),
	.combout(\Mux33~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~11 .lut_mask = 16'hEC64;
defparam \Mux33~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N19
dffeas \rfile[29][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][29] .is_wysiwyg = "true";
defparam \rfile[29][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N16
cycloneive_lcell_comb \rfile[25][29]~feeder (
// Equation(s):
// \rfile[25][29]~feeder_combout  = \wdat_WB[29]~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_29),
	.cin(gnd),
	.combout(\rfile[25][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[25][29]~feeder .lut_mask = 16'hFF00;
defparam \rfile[25][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N17
dffeas \rfile[25][29] (
	.clk(!CLK),
	.d(\rfile[25][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][29] .is_wysiwyg = "true";
defparam \rfile[25][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N21
dffeas \rfile[21][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][29] .is_wysiwyg = "true";
defparam \rfile[21][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N15
dffeas \rfile[17][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][29] .is_wysiwyg = "true";
defparam \rfile[17][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N20
cycloneive_lcell_comb \Mux34~0 (
// Equation(s):
// \Mux34~0_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[21][29]~q )))) # (!instruction_D[18] & (!instruction_D[19] & ((\rfile[17][29]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[21][29]~q ),
	.datad(\rfile[17][29]~q ),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~0 .lut_mask = 16'hB9A8;
defparam \Mux34~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N28
cycloneive_lcell_comb \Mux34~1 (
// Equation(s):
// \Mux34~1_combout  = (instruction_D[19] & ((\Mux34~0_combout  & (\rfile[29][29]~q )) # (!\Mux34~0_combout  & ((\rfile[25][29]~q ))))) # (!instruction_D[19] & (((\Mux34~0_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[29][29]~q ),
	.datac(\rfile[25][29]~q ),
	.datad(\Mux34~0_combout ),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~1 .lut_mask = 16'hDDA0;
defparam \Mux34~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N31
dffeas \rfile[20][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][29] .is_wysiwyg = "true";
defparam \rfile[20][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N8
cycloneive_lcell_comb \rfile[28][29]~feeder (
// Equation(s):
// \rfile[28][29]~feeder_combout  = \wdat_WB[29]~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_29),
	.cin(gnd),
	.combout(\rfile[28][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][29]~feeder .lut_mask = 16'hFF00;
defparam \rfile[28][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N9
dffeas \rfile[28][29] (
	.clk(!CLK),
	.d(\rfile[28][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][29] .is_wysiwyg = "true";
defparam \rfile[28][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N8
cycloneive_lcell_comb \Mux34~5 (
// Equation(s):
// \Mux34~5_combout  = (\Mux34~4_combout  & (((\rfile[28][29]~q )) # (!instruction_D[18]))) # (!\Mux34~4_combout  & (instruction_D[18] & (\rfile[20][29]~q )))

	.dataa(\Mux34~4_combout ),
	.datab(instruction_D_18),
	.datac(\rfile[20][29]~q ),
	.datad(\rfile[28][29]~q ),
	.cin(gnd),
	.combout(\Mux34~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~5 .lut_mask = 16'hEA62;
defparam \Mux34~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y36_N9
dffeas \rfile[30][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][29] .is_wysiwyg = "true";
defparam \rfile[30][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y35_N1
dffeas \rfile[22][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][29] .is_wysiwyg = "true";
defparam \rfile[22][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N2
cycloneive_lcell_comb \rfile[18][29]~feeder (
// Equation(s):
// \rfile[18][29]~feeder_combout  = \wdat_WB[29]~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_29),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[18][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[18][29]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[18][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N6
cycloneive_lcell_comb \Decoder0~10 (
// Equation(s):
// \Decoder0~10_combout  = (!wsel_WB[2] & (!wsel_WB[0] & \Decoder0~6_combout ))

	.dataa(wsel_WB_2),
	.datab(wsel_WB_0),
	.datac(gnd),
	.datad(\Decoder0~6_combout ),
	.cin(gnd),
	.combout(\Decoder0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~10 .lut_mask = 16'h1100;
defparam \Decoder0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y35_N3
dffeas \rfile[18][29] (
	.clk(!CLK),
	.d(\rfile[18][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][29] .is_wysiwyg = "true";
defparam \rfile[18][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N8
cycloneive_lcell_comb \rfile[26][29]~feeder (
// Equation(s):
// \rfile[26][29]~feeder_combout  = \wdat_WB[29]~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_29),
	.cin(gnd),
	.combout(\rfile[26][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[26][29]~feeder .lut_mask = 16'hFF00;
defparam \rfile[26][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y36_N9
dffeas \rfile[26][29] (
	.clk(!CLK),
	.d(\rfile[26][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][29] .is_wysiwyg = "true";
defparam \rfile[26][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N24
cycloneive_lcell_comb \Mux34~2 (
// Equation(s):
// \Mux34~2_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[26][29]~q )))) # (!instruction_D[19] & (!instruction_D[18] & (\rfile[18][29]~q )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][29]~q ),
	.datad(\rfile[26][29]~q ),
	.cin(gnd),
	.combout(\Mux34~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~2 .lut_mask = 16'hBA98;
defparam \Mux34~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N0
cycloneive_lcell_comb \Mux34~3 (
// Equation(s):
// \Mux34~3_combout  = (instruction_D[18] & ((\Mux34~2_combout  & (\rfile[30][29]~q )) # (!\Mux34~2_combout  & ((\rfile[22][29]~q ))))) # (!instruction_D[18] & (((\Mux34~2_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[30][29]~q ),
	.datac(\rfile[22][29]~q ),
	.datad(\Mux34~2_combout ),
	.cin(gnd),
	.combout(\Mux34~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~3 .lut_mask = 16'hDDA0;
defparam \Mux34~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N4
cycloneive_lcell_comb \Mux34~6 (
// Equation(s):
// \Mux34~6_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & ((\Mux34~3_combout ))) # (!instruction_D[17] & (\Mux34~5_combout ))))

	.dataa(instruction_D_16),
	.datab(\Mux34~5_combout ),
	.datac(\Mux34~3_combout ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux34~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~6 .lut_mask = 16'hFA44;
defparam \Mux34~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N27
dffeas \rfile[31][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][29] .is_wysiwyg = "true";
defparam \rfile[31][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N9
dffeas \rfile[23][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][29] .is_wysiwyg = "true";
defparam \rfile[23][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N7
dffeas \rfile[19][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][29] .is_wysiwyg = "true";
defparam \rfile[19][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N8
cycloneive_lcell_comb \Mux34~7 (
// Equation(s):
// \Mux34~7_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[23][29]~q )) # (!instruction_D[18] & ((\rfile[19][29]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[23][29]~q ),
	.datad(\rfile[19][29]~q ),
	.cin(gnd),
	.combout(\Mux34~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~7 .lut_mask = 16'hD9C8;
defparam \Mux34~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N1
dffeas \rfile[27][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][29] .is_wysiwyg = "true";
defparam \rfile[27][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N0
cycloneive_lcell_comb \Mux34~8 (
// Equation(s):
// \Mux34~8_combout  = (\Mux34~7_combout  & ((\rfile[31][29]~q ) # ((!instruction_D[19])))) # (!\Mux34~7_combout  & (((\rfile[27][29]~q  & instruction_D[19]))))

	.dataa(\rfile[31][29]~q ),
	.datab(\Mux34~7_combout ),
	.datac(\rfile[27][29]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux34~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~8 .lut_mask = 16'hB8CC;
defparam \Mux34~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N5
dffeas \rfile[11][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][29] .is_wysiwyg = "true";
defparam \rfile[11][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N21
dffeas \rfile[9][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][29] .is_wysiwyg = "true";
defparam \rfile[9][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N21
dffeas \rfile[10][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][29] .is_wysiwyg = "true";
defparam \rfile[10][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N11
dffeas \rfile[8][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][29] .is_wysiwyg = "true";
defparam \rfile[8][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N20
cycloneive_lcell_comb \Mux34~10 (
// Equation(s):
// \Mux34~10_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][29]~q )))) # (!instruction_D[17] & (!instruction_D[16] & ((\rfile[8][29]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[10][29]~q ),
	.datad(\rfile[8][29]~q ),
	.cin(gnd),
	.combout(\Mux34~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~10 .lut_mask = 16'hB9A8;
defparam \Mux34~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N20
cycloneive_lcell_comb \Mux34~11 (
// Equation(s):
// \Mux34~11_combout  = (instruction_D[16] & ((\Mux34~10_combout  & (\rfile[11][29]~q )) # (!\Mux34~10_combout  & ((\rfile[9][29]~q ))))) # (!instruction_D[16] & (((\Mux34~10_combout ))))

	.dataa(\rfile[11][29]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[9][29]~q ),
	.datad(\Mux34~10_combout ),
	.cin(gnd),
	.combout(\Mux34~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~11 .lut_mask = 16'hBBC0;
defparam \Mux34~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N15
dffeas \rfile[13][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][29] .is_wysiwyg = "true";
defparam \rfile[13][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N29
dffeas \rfile[12][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][29] .is_wysiwyg = "true";
defparam \rfile[12][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N28
cycloneive_lcell_comb \Mux34~17 (
// Equation(s):
// \Mux34~17_combout  = (instruction_D[17] & (((instruction_D[16])))) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[13][29]~q )) # (!instruction_D[16] & ((\rfile[12][29]~q )))))

	.dataa(instruction_D_17),
	.datab(\rfile[13][29]~q ),
	.datac(\rfile[12][29]~q ),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux34~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~17 .lut_mask = 16'hEE50;
defparam \Mux34~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N15
dffeas \rfile[15][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][29] .is_wysiwyg = "true";
defparam \rfile[15][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N29
dffeas \rfile[14][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][29] .is_wysiwyg = "true";
defparam \rfile[14][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N14
cycloneive_lcell_comb \Mux34~18 (
// Equation(s):
// \Mux34~18_combout  = (\Mux34~17_combout  & (((\rfile[15][29]~q )) # (!instruction_D[17]))) # (!\Mux34~17_combout  & (instruction_D[17] & ((\rfile[14][29]~q ))))

	.dataa(\Mux34~17_combout ),
	.datab(instruction_D_17),
	.datac(\rfile[15][29]~q ),
	.datad(\rfile[14][29]~q ),
	.cin(gnd),
	.combout(\Mux34~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~18 .lut_mask = 16'hE6A2;
defparam \Mux34~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N9
dffeas \rfile[6][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][29] .is_wysiwyg = "true";
defparam \rfile[6][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N20
cycloneive_lcell_comb \Decoder0~30 (
// Equation(s):
// \Decoder0~30_combout  = (wsel_WB[2] & (!wsel_WB[0] & \Decoder0~28_combout ))

	.dataa(wsel_WB_2),
	.datab(gnd),
	.datac(wsel_WB_0),
	.datad(\Decoder0~28_combout ),
	.cin(gnd),
	.combout(\Decoder0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~30 .lut_mask = 16'h0A00;
defparam \Decoder0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N7
dffeas \rfile[4][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][29] .is_wysiwyg = "true";
defparam \rfile[4][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N25
dffeas \rfile[5][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][29] .is_wysiwyg = "true";
defparam \rfile[5][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N6
cycloneive_lcell_comb \Mux34~12 (
// Equation(s):
// \Mux34~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][29]~q ))) # (!instruction_D[16] & (\rfile[4][29]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][29]~q ),
	.datad(\rfile[5][29]~q ),
	.cin(gnd),
	.combout(\Mux34~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~12 .lut_mask = 16'hDC98;
defparam \Mux34~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N8
cycloneive_lcell_comb \Mux34~13 (
// Equation(s):
// \Mux34~13_combout  = (instruction_D[17] & ((\Mux34~12_combout  & (\rfile[7][29]~q )) # (!\Mux34~12_combout  & ((\rfile[6][29]~q ))))) # (!instruction_D[17] & (((\Mux34~12_combout ))))

	.dataa(\rfile[7][29]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[6][29]~q ),
	.datad(\Mux34~12_combout ),
	.cin(gnd),
	.combout(\Mux34~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~13 .lut_mask = 16'hBBC0;
defparam \Mux34~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N31
dffeas \rfile[2][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][29] .is_wysiwyg = "true";
defparam \rfile[2][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y33_N21
dffeas \rfile[3][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][29] .is_wysiwyg = "true";
defparam \rfile[3][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N10
cycloneive_lcell_comb \rfile[1][29]~feeder (
// Equation(s):
// \rfile[1][29]~feeder_combout  = \wdat_WB[29]~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_29),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[1][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[1][29]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[1][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N11
dffeas \rfile[1][29] (
	.clk(!CLK),
	.d(\rfile[1][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][29] .is_wysiwyg = "true";
defparam \rfile[1][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N20
cycloneive_lcell_comb \Mux34~14 (
// Equation(s):
// \Mux34~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][29]~q )) # (!instruction_D[17] & ((\rfile[1][29]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[3][29]~q ),
	.datad(\rfile[1][29]~q ),
	.cin(gnd),
	.combout(\Mux34~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~14 .lut_mask = 16'hC480;
defparam \Mux34~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N30
cycloneive_lcell_comb \Mux34~15 (
// Equation(s):
// \Mux34~15_combout  = (\Mux34~14_combout ) # ((!instruction_D[16] & (instruction_D[17] & \rfile[2][29]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[2][29]~q ),
	.datad(\Mux34~14_combout ),
	.cin(gnd),
	.combout(\Mux34~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~15 .lut_mask = 16'hFF40;
defparam \Mux34~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N10
cycloneive_lcell_comb \Mux34~16 (
// Equation(s):
// \Mux34~16_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\Mux34~13_combout )) # (!instruction_D[18] & ((\Mux34~15_combout )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux34~13_combout ),
	.datad(\Mux34~15_combout ),
	.cin(gnd),
	.combout(\Mux34~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~16 .lut_mask = 16'hD9C8;
defparam \Mux34~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N11
dffeas \rfile[31][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][28] .is_wysiwyg = "true";
defparam \rfile[31][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N17
dffeas \rfile[23][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][28] .is_wysiwyg = "true";
defparam \rfile[23][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N1
dffeas \rfile[27][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][28] .is_wysiwyg = "true";
defparam \rfile[27][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N3
dffeas \rfile[19][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][28] .is_wysiwyg = "true";
defparam \rfile[19][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N0
cycloneive_lcell_comb \Mux35~7 (
// Equation(s):
// \Mux35~7_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[27][28]~q )) # (!instruction_D[19] & ((\rfile[19][28]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[27][28]~q ),
	.datad(\rfile[19][28]~q ),
	.cin(gnd),
	.combout(\Mux35~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~7 .lut_mask = 16'hD9C8;
defparam \Mux35~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N16
cycloneive_lcell_comb \Mux35~8 (
// Equation(s):
// \Mux35~8_combout  = (instruction_D[18] & ((\Mux35~7_combout  & (\rfile[31][28]~q )) # (!\Mux35~7_combout  & ((\rfile[23][28]~q ))))) # (!instruction_D[18] & (((\Mux35~7_combout ))))

	.dataa(\rfile[31][28]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[23][28]~q ),
	.datad(\Mux35~7_combout ),
	.cin(gnd),
	.combout(\Mux35~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~8 .lut_mask = 16'hBBC0;
defparam \Mux35~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N25
dffeas \rfile[24][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][28] .is_wysiwyg = "true";
defparam \rfile[24][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y31_N19
dffeas \rfile[16][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][28] .is_wysiwyg = "true";
defparam \rfile[16][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y31_N29
dffeas \rfile[20][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][28] .is_wysiwyg = "true";
defparam \rfile[20][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N18
cycloneive_lcell_comb \Mux35~4 (
// Equation(s):
// \Mux35~4_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[20][28]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[16][28]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[16][28]~q ),
	.datad(\rfile[20][28]~q ),
	.cin(gnd),
	.combout(\Mux35~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~4 .lut_mask = 16'hBA98;
defparam \Mux35~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N24
cycloneive_lcell_comb \Mux35~5 (
// Equation(s):
// \Mux35~5_combout  = (instruction_D[19] & ((\Mux35~4_combout  & (\rfile[28][28]~q )) # (!\Mux35~4_combout  & ((\rfile[24][28]~q ))))) # (!instruction_D[19] & (((\Mux35~4_combout ))))

	.dataa(\rfile[28][28]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[24][28]~q ),
	.datad(\Mux35~4_combout ),
	.cin(gnd),
	.combout(\Mux35~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~5 .lut_mask = 16'hBBC0;
defparam \Mux35~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y34_N21
dffeas \rfile[26][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][28] .is_wysiwyg = "true";
defparam \rfile[26][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y34_N23
dffeas \rfile[30][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][28] .is_wysiwyg = "true";
defparam \rfile[30][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y34_N7
dffeas \rfile[18][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][28] .is_wysiwyg = "true";
defparam \rfile[18][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y34_N17
dffeas \rfile[22][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][28] .is_wysiwyg = "true";
defparam \rfile[22][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N6
cycloneive_lcell_comb \Mux35~2 (
// Equation(s):
// \Mux35~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[22][28]~q ))) # (!instruction_D[18] & (\rfile[18][28]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][28]~q ),
	.datad(\rfile[22][28]~q ),
	.cin(gnd),
	.combout(\Mux35~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~2 .lut_mask = 16'hDC98;
defparam \Mux35~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N22
cycloneive_lcell_comb \Mux35~3 (
// Equation(s):
// \Mux35~3_combout  = (instruction_D[19] & ((\Mux35~2_combout  & ((\rfile[30][28]~q ))) # (!\Mux35~2_combout  & (\rfile[26][28]~q )))) # (!instruction_D[19] & (((\Mux35~2_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[26][28]~q ),
	.datac(\rfile[30][28]~q ),
	.datad(\Mux35~2_combout ),
	.cin(gnd),
	.combout(\Mux35~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~3 .lut_mask = 16'hF588;
defparam \Mux35~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N8
cycloneive_lcell_comb \Mux35~6 (
// Equation(s):
// \Mux35~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\Mux35~3_combout ))) # (!instruction_D[17] & (\Mux35~5_combout ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux35~5_combout ),
	.datad(\Mux35~3_combout ),
	.cin(gnd),
	.combout(\Mux35~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~6 .lut_mask = 16'hDC98;
defparam \Mux35~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N9
dffeas \rfile[21][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][28] .is_wysiwyg = "true";
defparam \rfile[21][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N11
dffeas \rfile[29][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][28] .is_wysiwyg = "true";
defparam \rfile[29][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N17
dffeas \rfile[17][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][28] .is_wysiwyg = "true";
defparam \rfile[17][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y30_N29
dffeas \rfile[25][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][28] .is_wysiwyg = "true";
defparam \rfile[25][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N16
cycloneive_lcell_comb \Mux35~0 (
// Equation(s):
// \Mux35~0_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[25][28]~q )))) # (!instruction_D[19] & (!instruction_D[18] & (\rfile[17][28]~q )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[17][28]~q ),
	.datad(\rfile[25][28]~q ),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~0 .lut_mask = 16'hBA98;
defparam \Mux35~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N10
cycloneive_lcell_comb \Mux35~1 (
// Equation(s):
// \Mux35~1_combout  = (instruction_D[18] & ((\Mux35~0_combout  & ((\rfile[29][28]~q ))) # (!\Mux35~0_combout  & (\rfile[21][28]~q )))) # (!instruction_D[18] & (((\Mux35~0_combout ))))

	.dataa(\rfile[21][28]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[29][28]~q ),
	.datad(\Mux35~0_combout ),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~1 .lut_mask = 16'hF388;
defparam \Mux35~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N8
cycloneive_lcell_comb \rfile[14][28]~feeder (
// Equation(s):
// \rfile[14][28]~feeder_combout  = \wdat_WB[28]~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_28),
	.cin(gnd),
	.combout(\rfile[14][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][28]~feeder .lut_mask = 16'hFF00;
defparam \rfile[14][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N9
dffeas \rfile[14][28] (
	.clk(!CLK),
	.d(\rfile[14][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][28] .is_wysiwyg = "true";
defparam \rfile[14][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N11
dffeas \rfile[15][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][28] .is_wysiwyg = "true";
defparam \rfile[15][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N19
dffeas \rfile[13][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][28] .is_wysiwyg = "true";
defparam \rfile[13][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N11
dffeas \rfile[12][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][28] .is_wysiwyg = "true";
defparam \rfile[12][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N18
cycloneive_lcell_comb \Mux35~17 (
// Equation(s):
// \Mux35~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][28]~q )))) # (!instruction_D[16] & (!instruction_D[17] & ((\rfile[12][28]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[13][28]~q ),
	.datad(\rfile[12][28]~q ),
	.cin(gnd),
	.combout(\Mux35~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~17 .lut_mask = 16'hB9A8;
defparam \Mux35~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N10
cycloneive_lcell_comb \Mux35~18 (
// Equation(s):
// \Mux35~18_combout  = (instruction_D[17] & ((\Mux35~17_combout  & ((\rfile[15][28]~q ))) # (!\Mux35~17_combout  & (\rfile[14][28]~q )))) # (!instruction_D[17] & (((\Mux35~17_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[14][28]~q ),
	.datac(\rfile[15][28]~q ),
	.datad(\Mux35~17_combout ),
	.cin(gnd),
	.combout(\Mux35~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~18 .lut_mask = 16'hF588;
defparam \Mux35~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N9
dffeas \rfile[3][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][28] .is_wysiwyg = "true";
defparam \rfile[3][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y33_N19
dffeas \rfile[1][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][28] .is_wysiwyg = "true";
defparam \rfile[1][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N8
cycloneive_lcell_comb \Mux35~14 (
// Equation(s):
// \Mux35~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][28]~q )) # (!instruction_D[17] & ((\rfile[1][28]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[3][28]~q ),
	.datad(\rfile[1][28]~q ),
	.cin(gnd),
	.combout(\Mux35~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~14 .lut_mask = 16'hC480;
defparam \Mux35~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y33_N23
dffeas \rfile[2][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][28] .is_wysiwyg = "true";
defparam \rfile[2][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N16
cycloneive_lcell_comb \Mux35~15 (
// Equation(s):
// \Mux35~15_combout  = (\Mux35~14_combout ) # ((instruction_D[17] & (!instruction_D[16] & \rfile[2][28]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux35~14_combout ),
	.datad(\rfile[2][28]~q ),
	.cin(gnd),
	.combout(\Mux35~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~15 .lut_mask = 16'hF2F0;
defparam \Mux35~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N24
cycloneive_lcell_comb \rfile[11][28]~feeder (
// Equation(s):
// \rfile[11][28]~feeder_combout  = \wdat_WB[28]~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_28),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[11][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][28]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[11][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y33_N25
dffeas \rfile[11][28] (
	.clk(!CLK),
	.d(\rfile[11][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][28] .is_wysiwyg = "true";
defparam \rfile[11][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N11
dffeas \rfile[9][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][28] .is_wysiwyg = "true";
defparam \rfile[9][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N19
dffeas \rfile[8][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][28] .is_wysiwyg = "true";
defparam \rfile[8][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N13
dffeas \rfile[10][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][28] .is_wysiwyg = "true";
defparam \rfile[10][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N18
cycloneive_lcell_comb \Mux35~12 (
// Equation(s):
// \Mux35~12_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][28]~q )))) # (!instruction_D[17] & (!instruction_D[16] & (\rfile[8][28]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[8][28]~q ),
	.datad(\rfile[10][28]~q ),
	.cin(gnd),
	.combout(\Mux35~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~12 .lut_mask = 16'hBA98;
defparam \Mux35~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N10
cycloneive_lcell_comb \Mux35~13 (
// Equation(s):
// \Mux35~13_combout  = (instruction_D[16] & ((\Mux35~12_combout  & (\rfile[11][28]~q )) # (!\Mux35~12_combout  & ((\rfile[9][28]~q ))))) # (!instruction_D[16] & (((\Mux35~12_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][28]~q ),
	.datac(\rfile[9][28]~q ),
	.datad(\Mux35~12_combout ),
	.cin(gnd),
	.combout(\Mux35~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~13 .lut_mask = 16'hDDA0;
defparam \Mux35~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N16
cycloneive_lcell_comb \Mux35~16 (
// Equation(s):
// \Mux35~16_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\Mux35~13_combout ))) # (!instruction_D[19] & (\Mux35~15_combout ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\Mux35~15_combout ),
	.datad(\Mux35~13_combout ),
	.cin(gnd),
	.combout(\Mux35~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~16 .lut_mask = 16'hDC98;
defparam \Mux35~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N15
dffeas \rfile[4][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][28] .is_wysiwyg = "true";
defparam \rfile[4][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N21
dffeas \rfile[5][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][28] .is_wysiwyg = "true";
defparam \rfile[5][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N14
cycloneive_lcell_comb \Mux35~10 (
// Equation(s):
// \Mux35~10_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][28]~q ))) # (!instruction_D[16] & (\rfile[4][28]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][28]~q ),
	.datad(\rfile[5][28]~q ),
	.cin(gnd),
	.combout(\Mux35~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~10 .lut_mask = 16'hDC98;
defparam \Mux35~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N7
dffeas \rfile[7][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][28] .is_wysiwyg = "true";
defparam \rfile[7][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y36_N21
dffeas \rfile[6][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][28] .is_wysiwyg = "true";
defparam \rfile[6][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N6
cycloneive_lcell_comb \Mux35~11 (
// Equation(s):
// \Mux35~11_combout  = (instruction_D[17] & ((\Mux35~10_combout  & (\rfile[7][28]~q )) # (!\Mux35~10_combout  & ((\rfile[6][28]~q ))))) # (!instruction_D[17] & (\Mux35~10_combout ))

	.dataa(instruction_D_17),
	.datab(\Mux35~10_combout ),
	.datac(\rfile[7][28]~q ),
	.datad(\rfile[6][28]~q ),
	.cin(gnd),
	.combout(\Mux35~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~11 .lut_mask = 16'hE6C4;
defparam \Mux35~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N19
dffeas \rfile[31][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][27] .is_wysiwyg = "true";
defparam \rfile[31][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y29_N29
dffeas \rfile[27][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][27] .is_wysiwyg = "true";
defparam \rfile[27][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N29
dffeas \rfile[23][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][27] .is_wysiwyg = "true";
defparam \rfile[23][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N28
cycloneive_lcell_comb \Mux36~7 (
// Equation(s):
// \Mux36~7_combout  = (instruction_D[18] & (((\rfile[23][27]~q ) # (instruction_D[19])))) # (!instruction_D[18] & (\rfile[19][27]~q  & ((!instruction_D[19]))))

	.dataa(\rfile[19][27]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[23][27]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux36~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~7 .lut_mask = 16'hCCE2;
defparam \Mux36~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N28
cycloneive_lcell_comb \Mux36~8 (
// Equation(s):
// \Mux36~8_combout  = (instruction_D[19] & ((\Mux36~7_combout  & (\rfile[31][27]~q )) # (!\Mux36~7_combout  & ((\rfile[27][27]~q ))))) # (!instruction_D[19] & (((\Mux36~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[31][27]~q ),
	.datac(\rfile[27][27]~q ),
	.datad(\Mux36~7_combout ),
	.cin(gnd),
	.combout(\Mux36~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~8 .lut_mask = 16'hDDA0;
defparam \Mux36~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N10
cycloneive_lcell_comb \rfile[25][27]~feeder (
// Equation(s):
// \rfile[25][27]~feeder_combout  = \wdat_WB[27]~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_27),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[25][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[25][27]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[25][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N11
dffeas \rfile[25][27] (
	.clk(!CLK),
	.d(\rfile[25][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][27] .is_wysiwyg = "true";
defparam \rfile[25][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N1
dffeas \rfile[29][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][27] .is_wysiwyg = "true";
defparam \rfile[29][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N23
dffeas \rfile[17][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][27] .is_wysiwyg = "true";
defparam \rfile[17][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N9
dffeas \rfile[21][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][27] .is_wysiwyg = "true";
defparam \rfile[21][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N22
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[21][27]~q ))) # (!instruction_D[18] & (\rfile[17][27]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[17][27]~q ),
	.datad(\rfile[21][27]~q ),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'hDC98;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N0
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (instruction_D[19] & ((\Mux36~0_combout  & ((\rfile[29][27]~q ))) # (!\Mux36~0_combout  & (\rfile[25][27]~q )))) # (!instruction_D[19] & (((\Mux36~0_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[25][27]~q ),
	.datac(\rfile[29][27]~q ),
	.datad(\Mux36~0_combout ),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'hF588;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y36_N13
dffeas \rfile[30][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][27] .is_wysiwyg = "true";
defparam \rfile[30][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y36_N3
dffeas \rfile[26][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][27] .is_wysiwyg = "true";
defparam \rfile[26][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y36_N19
dffeas \rfile[18][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][27] .is_wysiwyg = "true";
defparam \rfile[18][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N2
cycloneive_lcell_comb \Mux36~2 (
// Equation(s):
// \Mux36~2_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[26][27]~q )) # (!instruction_D[19] & ((\rfile[18][27]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[26][27]~q ),
	.datad(\rfile[18][27]~q ),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~2 .lut_mask = 16'hD9C8;
defparam \Mux36~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N12
cycloneive_lcell_comb \Mux36~3 (
// Equation(s):
// \Mux36~3_combout  = (instruction_D[18] & ((\Mux36~2_combout  & ((\rfile[30][27]~q ))) # (!\Mux36~2_combout  & (\rfile[22][27]~q )))) # (!instruction_D[18] & (((\Mux36~2_combout ))))

	.dataa(\rfile[22][27]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[30][27]~q ),
	.datad(\Mux36~2_combout ),
	.cin(gnd),
	.combout(\Mux36~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~3 .lut_mask = 16'hF388;
defparam \Mux36~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y32_N19
dffeas \rfile[24][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][27] .is_wysiwyg = "true";
defparam \rfile[24][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N17
dffeas \rfile[16][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][27] .is_wysiwyg = "true";
defparam \rfile[16][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N18
cycloneive_lcell_comb \Mux36~4 (
// Equation(s):
// \Mux36~4_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[24][27]~q )) # (!instruction_D[19] & ((\rfile[16][27]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[24][27]~q ),
	.datad(\rfile[16][27]~q ),
	.cin(gnd),
	.combout(\Mux36~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~4 .lut_mask = 16'hD9C8;
defparam \Mux36~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N22
cycloneive_lcell_comb \rfile[20][27]~feeder (
// Equation(s):
// \rfile[20][27]~feeder_combout  = \wdat_WB[27]~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_27),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[20][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[20][27]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[20][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N23
dffeas \rfile[20][27] (
	.clk(!CLK),
	.d(\rfile[20][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][27] .is_wysiwyg = "true";
defparam \rfile[20][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N0
cycloneive_lcell_comb \Mux36~5 (
// Equation(s):
// \Mux36~5_combout  = (instruction_D[18] & ((\Mux36~4_combout  & (\rfile[28][27]~q )) # (!\Mux36~4_combout  & ((\rfile[20][27]~q ))))) # (!instruction_D[18] & (((\Mux36~4_combout ))))

	.dataa(\rfile[28][27]~q ),
	.datab(instruction_D_18),
	.datac(\Mux36~4_combout ),
	.datad(\rfile[20][27]~q ),
	.cin(gnd),
	.combout(\Mux36~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~5 .lut_mask = 16'hBCB0;
defparam \Mux36~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N26
cycloneive_lcell_comb \Mux36~6 (
// Equation(s):
// \Mux36~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux36~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & ((\Mux36~5_combout ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux36~3_combout ),
	.datad(\Mux36~5_combout ),
	.cin(gnd),
	.combout(\Mux36~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~6 .lut_mask = 16'hB9A8;
defparam \Mux36~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N13
dffeas \rfile[13][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][27] .is_wysiwyg = "true";
defparam \rfile[13][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N7
dffeas \rfile[12][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][27] .is_wysiwyg = "true";
defparam \rfile[12][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N12
cycloneive_lcell_comb \Mux36~17 (
// Equation(s):
// \Mux36~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][27]~q )))) # (!instruction_D[16] & (!instruction_D[17] & ((\rfile[12][27]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[13][27]~q ),
	.datad(\rfile[12][27]~q ),
	.cin(gnd),
	.combout(\Mux36~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~17 .lut_mask = 16'hB9A8;
defparam \Mux36~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N23
dffeas \rfile[14][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][27] .is_wysiwyg = "true";
defparam \rfile[14][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N17
dffeas \rfile[15][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][27] .is_wysiwyg = "true";
defparam \rfile[15][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N22
cycloneive_lcell_comb \Mux36~18 (
// Equation(s):
// \Mux36~18_combout  = (\Mux36~17_combout  & (((\rfile[15][27]~q )) # (!instruction_D[17]))) # (!\Mux36~17_combout  & (instruction_D[17] & (\rfile[14][27]~q )))

	.dataa(\Mux36~17_combout ),
	.datab(instruction_D_17),
	.datac(\rfile[14][27]~q ),
	.datad(\rfile[15][27]~q ),
	.cin(gnd),
	.combout(\Mux36~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~18 .lut_mask = 16'hEA62;
defparam \Mux36~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N29
dffeas \rfile[6][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][27] .is_wysiwyg = "true";
defparam \rfile[6][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N29
dffeas \rfile[5][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][27] .is_wysiwyg = "true";
defparam \rfile[5][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N11
dffeas \rfile[4][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][27] .is_wysiwyg = "true";
defparam \rfile[4][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N28
cycloneive_lcell_comb \Mux36~12 (
// Equation(s):
// \Mux36~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[5][27]~q )) # (!instruction_D[16] & ((\rfile[4][27]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[5][27]~q ),
	.datad(\rfile[4][27]~q ),
	.cin(gnd),
	.combout(\Mux36~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~12 .lut_mask = 16'hD9C8;
defparam \Mux36~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N28
cycloneive_lcell_comb \Mux36~13 (
// Equation(s):
// \Mux36~13_combout  = (instruction_D[17] & ((\Mux36~12_combout  & (\rfile[7][27]~q )) # (!\Mux36~12_combout  & ((\rfile[6][27]~q ))))) # (!instruction_D[17] & (((\Mux36~12_combout ))))

	.dataa(\rfile[7][27]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[6][27]~q ),
	.datad(\Mux36~12_combout ),
	.cin(gnd),
	.combout(\Mux36~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~13 .lut_mask = 16'hBBC0;
defparam \Mux36~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y33_N21
dffeas \rfile[2][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][27] .is_wysiwyg = "true";
defparam \rfile[2][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y33_N23
dffeas \rfile[1][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][27] .is_wysiwyg = "true";
defparam \rfile[1][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N3
dffeas \rfile[3][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][27] .is_wysiwyg = "true";
defparam \rfile[3][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N18
cycloneive_lcell_comb \Mux36~14 (
// Equation(s):
// \Mux36~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][27]~q ))) # (!instruction_D[17] & (\rfile[1][27]~q ))))

	.dataa(instruction_D_17),
	.datab(\rfile[1][27]~q ),
	.datac(instruction_D_16),
	.datad(\rfile[3][27]~q ),
	.cin(gnd),
	.combout(\Mux36~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~14 .lut_mask = 16'hE040;
defparam \Mux36~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N20
cycloneive_lcell_comb \Mux36~15 (
// Equation(s):
// \Mux36~15_combout  = (\Mux36~14_combout ) # ((instruction_D[17] & (!instruction_D[16] & \rfile[2][27]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[2][27]~q ),
	.datad(\Mux36~14_combout ),
	.cin(gnd),
	.combout(\Mux36~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~15 .lut_mask = 16'hFF20;
defparam \Mux36~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N14
cycloneive_lcell_comb \Mux36~16 (
// Equation(s):
// \Mux36~16_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\Mux36~13_combout )) # (!instruction_D[18] & ((\Mux36~15_combout )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux36~13_combout ),
	.datad(\Mux36~15_combout ),
	.cin(gnd),
	.combout(\Mux36~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~16 .lut_mask = 16'hD9C8;
defparam \Mux36~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N10
cycloneive_lcell_comb \rfile[11][27]~feeder (
// Equation(s):
// \rfile[11][27]~feeder_combout  = \wdat_WB[27]~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_27),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[11][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][27]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[11][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y33_N11
dffeas \rfile[11][27] (
	.clk(!CLK),
	.d(\rfile[11][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][27] .is_wysiwyg = "true";
defparam \rfile[11][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N31
dffeas \rfile[8][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][27] .is_wysiwyg = "true";
defparam \rfile[8][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N17
dffeas \rfile[10][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][27] .is_wysiwyg = "true";
defparam \rfile[10][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N30
cycloneive_lcell_comb \Mux36~10 (
// Equation(s):
// \Mux36~10_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][27]~q )))) # (!instruction_D[17] & (!instruction_D[16] & (\rfile[8][27]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[8][27]~q ),
	.datad(\rfile[10][27]~q ),
	.cin(gnd),
	.combout(\Mux36~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~10 .lut_mask = 16'hBA98;
defparam \Mux36~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N21
dffeas \rfile[9][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][27] .is_wysiwyg = "true";
defparam \rfile[9][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N28
cycloneive_lcell_comb \Mux36~11 (
// Equation(s):
// \Mux36~11_combout  = (instruction_D[16] & ((\Mux36~10_combout  & (\rfile[11][27]~q )) # (!\Mux36~10_combout  & ((\rfile[9][27]~q ))))) # (!instruction_D[16] & (((\Mux36~10_combout ))))

	.dataa(\rfile[11][27]~q ),
	.datab(instruction_D_16),
	.datac(\Mux36~10_combout ),
	.datad(\rfile[9][27]~q ),
	.cin(gnd),
	.combout(\Mux36~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~11 .lut_mask = 16'hBCB0;
defparam \Mux36~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N22
cycloneive_lcell_comb \rfile[31][26]~feeder (
// Equation(s):
// \rfile[31][26]~feeder_combout  = \wdat_WB[26]~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_26),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[31][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[31][26]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[31][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N23
dffeas \rfile[31][26] (
	.clk(!CLK),
	.d(\rfile[31][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][26] .is_wysiwyg = "true";
defparam \rfile[31][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N25
dffeas \rfile[23][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][26] .is_wysiwyg = "true";
defparam \rfile[23][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N17
dffeas \rfile[27][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][26] .is_wysiwyg = "true";
defparam \rfile[27][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N11
dffeas \rfile[19][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][26] .is_wysiwyg = "true";
defparam \rfile[19][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N16
cycloneive_lcell_comb \Mux37~7 (
// Equation(s):
// \Mux37~7_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[27][26]~q )) # (!instruction_D[19] & ((\rfile[19][26]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[27][26]~q ),
	.datad(\rfile[19][26]~q ),
	.cin(gnd),
	.combout(\Mux37~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~7 .lut_mask = 16'hD9C8;
defparam \Mux37~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N24
cycloneive_lcell_comb \Mux37~8 (
// Equation(s):
// \Mux37~8_combout  = (instruction_D[18] & ((\Mux37~7_combout  & (\rfile[31][26]~q )) # (!\Mux37~7_combout  & ((\rfile[23][26]~q ))))) # (!instruction_D[18] & (((\Mux37~7_combout ))))

	.dataa(\rfile[31][26]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[23][26]~q ),
	.datad(\Mux37~7_combout ),
	.cin(gnd),
	.combout(\Mux37~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~8 .lut_mask = 16'hBBC0;
defparam \Mux37~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N1
dffeas \rfile[24][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][26] .is_wysiwyg = "true";
defparam \rfile[24][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N7
dffeas \rfile[28][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][26] .is_wysiwyg = "true";
defparam \rfile[28][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N0
cycloneive_lcell_comb \Mux37~5 (
// Equation(s):
// \Mux37~5_combout  = (\Mux37~4_combout  & (((\rfile[28][26]~q )) # (!instruction_D[19]))) # (!\Mux37~4_combout  & (instruction_D[19] & (\rfile[24][26]~q )))

	.dataa(\Mux37~4_combout ),
	.datab(instruction_D_19),
	.datac(\rfile[24][26]~q ),
	.datad(\rfile[28][26]~q ),
	.cin(gnd),
	.combout(\Mux37~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~5 .lut_mask = 16'hEA62;
defparam \Mux37~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y34_N9
dffeas \rfile[22][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][26] .is_wysiwyg = "true";
defparam \rfile[22][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N8
cycloneive_lcell_comb \Mux37~2 (
// Equation(s):
// \Mux37~2_combout  = (instruction_D[18] & (((\rfile[22][26]~q ) # (instruction_D[19])))) # (!instruction_D[18] & (\rfile[18][26]~q  & ((!instruction_D[19]))))

	.dataa(\rfile[18][26]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[22][26]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux37~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~2 .lut_mask = 16'hCCE2;
defparam \Mux37~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y34_N13
dffeas \rfile[26][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][26] .is_wysiwyg = "true";
defparam \rfile[26][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N1
dffeas \rfile[30][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][26] .is_wysiwyg = "true";
defparam \rfile[30][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N12
cycloneive_lcell_comb \Mux37~3 (
// Equation(s):
// \Mux37~3_combout  = (instruction_D[19] & ((\Mux37~2_combout  & ((\rfile[30][26]~q ))) # (!\Mux37~2_combout  & (\rfile[26][26]~q )))) # (!instruction_D[19] & (\Mux37~2_combout ))

	.dataa(instruction_D_19),
	.datab(\Mux37~2_combout ),
	.datac(\rfile[26][26]~q ),
	.datad(\rfile[30][26]~q ),
	.cin(gnd),
	.combout(\Mux37~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~3 .lut_mask = 16'hEC64;
defparam \Mux37~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N22
cycloneive_lcell_comb \Mux37~6 (
// Equation(s):
// \Mux37~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux37~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & (\Mux37~5_combout )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux37~5_combout ),
	.datad(\Mux37~3_combout ),
	.cin(gnd),
	.combout(\Mux37~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~6 .lut_mask = 16'hBA98;
defparam \Mux37~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N16
cycloneive_lcell_comb \rfile[29][26]~feeder (
// Equation(s):
// \rfile[29][26]~feeder_combout  = \wdat_WB[26]~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_26),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[29][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[29][26]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[29][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N17
dffeas \rfile[29][26] (
	.clk(!CLK),
	.d(\rfile[29][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][26] .is_wysiwyg = "true";
defparam \rfile[29][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N22
cycloneive_lcell_comb \rfile[21][26]~feeder (
// Equation(s):
// \rfile[21][26]~feeder_combout  = \wdat_WB[26]~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_26),
	.cin(gnd),
	.combout(\rfile[21][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][26]~feeder .lut_mask = 16'hFF00;
defparam \rfile[21][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N23
dffeas \rfile[21][26] (
	.clk(!CLK),
	.d(\rfile[21][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][26] .is_wysiwyg = "true";
defparam \rfile[21][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N29
dffeas \rfile[25][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][26] .is_wysiwyg = "true";
defparam \rfile[25][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N28
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[25][26]~q ))) # (!instruction_D[19] & (\rfile[17][26]~q ))))

	.dataa(\rfile[17][26]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[25][26]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hFC22;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N22
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (instruction_D[18] & ((\Mux37~0_combout  & (\rfile[29][26]~q )) # (!\Mux37~0_combout  & ((\rfile[21][26]~q ))))) # (!instruction_D[18] & (((\Mux37~0_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[29][26]~q ),
	.datac(\rfile[21][26]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hDDA0;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N10
cycloneive_lcell_comb \rfile[9][26]~feeder (
// Equation(s):
// \rfile[9][26]~feeder_combout  = \wdat_WB[26]~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_26),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[9][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][26]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[9][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N11
dffeas \rfile[9][26] (
	.clk(!CLK),
	.d(\rfile[9][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][26] .is_wysiwyg = "true";
defparam \rfile[9][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N7
dffeas \rfile[8][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][26] .is_wysiwyg = "true";
defparam \rfile[8][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N6
cycloneive_lcell_comb \Mux37~12 (
// Equation(s):
// \Mux37~12_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & (\rfile[10][26]~q )) # (!instruction_D[17] & ((\rfile[8][26]~q )))))

	.dataa(\rfile[10][26]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[8][26]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux37~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~12 .lut_mask = 16'hEE30;
defparam \Mux37~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N30
cycloneive_lcell_comb \Mux37~13 (
// Equation(s):
// \Mux37~13_combout  = (instruction_D[16] & ((\Mux37~12_combout  & (\rfile[11][26]~q )) # (!\Mux37~12_combout  & ((\rfile[9][26]~q ))))) # (!instruction_D[16] & (((\Mux37~12_combout ))))

	.dataa(\rfile[11][26]~q ),
	.datab(\rfile[9][26]~q ),
	.datac(instruction_D_16),
	.datad(\Mux37~12_combout ),
	.cin(gnd),
	.combout(\Mux37~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~13 .lut_mask = 16'hAFC0;
defparam \Mux37~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N10
cycloneive_lcell_comb \rfile[2][26]~feeder (
// Equation(s):
// \rfile[2][26]~feeder_combout  = \wdat_WB[26]~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_26),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[2][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][26]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[2][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N11
dffeas \rfile[2][26] (
	.clk(!CLK),
	.d(\rfile[2][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][26] .is_wysiwyg = "true";
defparam \rfile[2][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N25
dffeas \rfile[3][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][26] .is_wysiwyg = "true";
defparam \rfile[3][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N7
dffeas \rfile[1][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][26] .is_wysiwyg = "true";
defparam \rfile[1][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N6
cycloneive_lcell_comb \Mux37~14 (
// Equation(s):
// \Mux37~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][26]~q )) # (!instruction_D[17] & ((\rfile[1][26]~q )))))

	.dataa(instruction_D_16),
	.datab(\rfile[3][26]~q ),
	.datac(\rfile[1][26]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux37~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~14 .lut_mask = 16'h88A0;
defparam \Mux37~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N12
cycloneive_lcell_comb \Mux37~15 (
// Equation(s):
// \Mux37~15_combout  = (\Mux37~14_combout ) # ((instruction_D[17] & (\rfile[2][26]~q  & !instruction_D[16])))

	.dataa(instruction_D_17),
	.datab(\rfile[2][26]~q ),
	.datac(instruction_D_16),
	.datad(\Mux37~14_combout ),
	.cin(gnd),
	.combout(\Mux37~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~15 .lut_mask = 16'hFF08;
defparam \Mux37~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N10
cycloneive_lcell_comb \Mux37~16 (
// Equation(s):
// \Mux37~16_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\Mux37~13_combout )) # (!instruction_D[19] & ((\Mux37~15_combout )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\Mux37~13_combout ),
	.datad(\Mux37~15_combout ),
	.cin(gnd),
	.combout(\Mux37~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~16 .lut_mask = 16'hD9C8;
defparam \Mux37~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N19
dffeas \rfile[4][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][26] .is_wysiwyg = "true";
defparam \rfile[4][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N17
dffeas \rfile[5][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][26] .is_wysiwyg = "true";
defparam \rfile[5][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N18
cycloneive_lcell_comb \Mux37~10 (
// Equation(s):
// \Mux37~10_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][26]~q ))) # (!instruction_D[16] & (\rfile[4][26]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][26]~q ),
	.datad(\rfile[5][26]~q ),
	.cin(gnd),
	.combout(\Mux37~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~10 .lut_mask = 16'hDC98;
defparam \Mux37~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N19
dffeas \rfile[7][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][26] .is_wysiwyg = "true";
defparam \rfile[7][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y36_N13
dffeas \rfile[6][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][26] .is_wysiwyg = "true";
defparam \rfile[6][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N18
cycloneive_lcell_comb \Mux37~11 (
// Equation(s):
// \Mux37~11_combout  = (instruction_D[17] & ((\Mux37~10_combout  & (\rfile[7][26]~q )) # (!\Mux37~10_combout  & ((\rfile[6][26]~q ))))) # (!instruction_D[17] & (\Mux37~10_combout ))

	.dataa(instruction_D_17),
	.datab(\Mux37~10_combout ),
	.datac(\rfile[7][26]~q ),
	.datad(\rfile[6][26]~q ),
	.cin(gnd),
	.combout(\Mux37~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~11 .lut_mask = 16'hE6C4;
defparam \Mux37~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N11
dffeas \rfile[12][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][26] .is_wysiwyg = "true";
defparam \rfile[12][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N21
dffeas \rfile[13][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][26] .is_wysiwyg = "true";
defparam \rfile[13][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N10
cycloneive_lcell_comb \Mux37~17 (
// Equation(s):
// \Mux37~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][26]~q )))) # (!instruction_D[16] & (!instruction_D[17] & (\rfile[12][26]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[12][26]~q ),
	.datad(\rfile[13][26]~q ),
	.cin(gnd),
	.combout(\Mux37~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~17 .lut_mask = 16'hBA98;
defparam \Mux37~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N7
dffeas \rfile[14][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][26] .is_wysiwyg = "true";
defparam \rfile[14][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N25
dffeas \rfile[15][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][26] .is_wysiwyg = "true";
defparam \rfile[15][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N6
cycloneive_lcell_comb \Mux37~18 (
// Equation(s):
// \Mux37~18_combout  = (\Mux37~17_combout  & (((\rfile[15][26]~q )) # (!instruction_D[17]))) # (!\Mux37~17_combout  & (instruction_D[17] & (\rfile[14][26]~q )))

	.dataa(\Mux37~17_combout ),
	.datab(instruction_D_17),
	.datac(\rfile[14][26]~q ),
	.datad(\rfile[15][26]~q ),
	.cin(gnd),
	.combout(\Mux37~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~18 .lut_mask = 16'hEA62;
defparam \Mux37~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y29_N25
dffeas \rfile[23][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][25] .is_wysiwyg = "true";
defparam \rfile[23][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N24
cycloneive_lcell_comb \Mux38~7 (
// Equation(s):
// \Mux38~7_combout  = (instruction_D[18] & (((\rfile[23][25]~q ) # (instruction_D[19])))) # (!instruction_D[18] & (\rfile[19][25]~q  & ((!instruction_D[19]))))

	.dataa(\rfile[19][25]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[23][25]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux38~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~7 .lut_mask = 16'hCCE2;
defparam \Mux38~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N15
dffeas \rfile[31][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][25] .is_wysiwyg = "true";
defparam \rfile[31][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y29_N21
dffeas \rfile[27][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][25] .is_wysiwyg = "true";
defparam \rfile[27][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N20
cycloneive_lcell_comb \Mux38~8 (
// Equation(s):
// \Mux38~8_combout  = (\Mux38~7_combout  & ((\rfile[31][25]~q ) # ((!instruction_D[19])))) # (!\Mux38~7_combout  & (((\rfile[27][25]~q  & instruction_D[19]))))

	.dataa(\Mux38~7_combout ),
	.datab(\rfile[31][25]~q ),
	.datac(\rfile[27][25]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux38~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~8 .lut_mask = 16'hD8AA;
defparam \Mux38~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N15
dffeas \rfile[29][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][25] .is_wysiwyg = "true";
defparam \rfile[29][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N29
dffeas \rfile[25][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][25] .is_wysiwyg = "true";
defparam \rfile[25][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N1
dffeas \rfile[17][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][25] .is_wysiwyg = "true";
defparam \rfile[17][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N20
cycloneive_lcell_comb \rfile[21][25]~feeder (
// Equation(s):
// \rfile[21][25]~feeder_combout  = \wdat_WB[25]~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_25),
	.cin(gnd),
	.combout(\rfile[21][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][25]~feeder .lut_mask = 16'hFF00;
defparam \rfile[21][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N21
dffeas \rfile[21][25] (
	.clk(!CLK),
	.d(\rfile[21][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][25] .is_wysiwyg = "true";
defparam \rfile[21][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N2
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[21][25]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[17][25]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[17][25]~q ),
	.datad(\rfile[21][25]~q ),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hBA98;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N28
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (instruction_D[19] & ((\Mux38~0_combout  & (\rfile[29][25]~q )) # (!\Mux38~0_combout  & ((\rfile[25][25]~q ))))) # (!instruction_D[19] & (((\Mux38~0_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[29][25]~q ),
	.datac(\rfile[25][25]~q ),
	.datad(\Mux38~0_combout ),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hDDA0;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N9
dffeas \rfile[22][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][25] .is_wysiwyg = "true";
defparam \rfile[22][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N18
cycloneive_lcell_comb \rfile[30][25]~feeder (
// Equation(s):
// \rfile[30][25]~feeder_combout  = \wdat_WB[25]~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[30][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[30][25]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[30][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N19
dffeas \rfile[30][25] (
	.clk(!CLK),
	.d(\rfile[30][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][25] .is_wysiwyg = "true";
defparam \rfile[30][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N8
cycloneive_lcell_comb \Mux38~3 (
// Equation(s):
// \Mux38~3_combout  = (\Mux38~2_combout  & (((\rfile[30][25]~q )) # (!instruction_D[18]))) # (!\Mux38~2_combout  & (instruction_D[18] & (\rfile[22][25]~q )))

	.dataa(\Mux38~2_combout ),
	.datab(instruction_D_18),
	.datac(\rfile[22][25]~q ),
	.datad(\rfile[30][25]~q ),
	.cin(gnd),
	.combout(\Mux38~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~3 .lut_mask = 16'hEA62;
defparam \Mux38~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y31_N13
dffeas \rfile[20][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][25] .is_wysiwyg = "true";
defparam \rfile[20][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y31_N3
dffeas \rfile[16][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][25] .is_wysiwyg = "true";
defparam \rfile[16][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X77_Y32_N28
cycloneive_lcell_comb \rfile[24][25]~feeder (
// Equation(s):
// \rfile[24][25]~feeder_combout  = \wdat_WB[25]~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[24][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[24][25]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[24][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X77_Y32_N29
dffeas \rfile[24][25] (
	.clk(!CLK),
	.d(\rfile[24][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][25] .is_wysiwyg = "true";
defparam \rfile[24][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N2
cycloneive_lcell_comb \Mux38~4 (
// Equation(s):
// \Mux38~4_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[24][25]~q ))) # (!instruction_D[19] & (\rfile[16][25]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[16][25]~q ),
	.datad(\rfile[24][25]~q ),
	.cin(gnd),
	.combout(\Mux38~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~4 .lut_mask = 16'hDC98;
defparam \Mux38~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N12
cycloneive_lcell_comb \Mux38~5 (
// Equation(s):
// \Mux38~5_combout  = (instruction_D[18] & ((\Mux38~4_combout  & (\rfile[28][25]~q )) # (!\Mux38~4_combout  & ((\rfile[20][25]~q ))))) # (!instruction_D[18] & (((\Mux38~4_combout ))))

	.dataa(\rfile[28][25]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[20][25]~q ),
	.datad(\Mux38~4_combout ),
	.cin(gnd),
	.combout(\Mux38~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~5 .lut_mask = 16'hBBC0;
defparam \Mux38~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N12
cycloneive_lcell_comb \Mux38~6 (
// Equation(s):
// \Mux38~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\Mux38~3_combout )) # (!instruction_D[17] & ((\Mux38~5_combout )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux38~3_combout ),
	.datad(\Mux38~5_combout ),
	.cin(gnd),
	.combout(\Mux38~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~6 .lut_mask = 16'hD9C8;
defparam \Mux38~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N5
dffeas \rfile[14][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][25] .is_wysiwyg = "true";
defparam \rfile[14][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N31
dffeas \rfile[15][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][25] .is_wysiwyg = "true";
defparam \rfile[15][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N13
dffeas \rfile[12][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][25] .is_wysiwyg = "true";
defparam \rfile[12][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N17
dffeas \rfile[13][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][25] .is_wysiwyg = "true";
defparam \rfile[13][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N12
cycloneive_lcell_comb \Mux38~17 (
// Equation(s):
// \Mux38~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][25]~q ))) # (!instruction_D[16] & (\rfile[12][25]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][25]~q ),
	.datad(\rfile[13][25]~q ),
	.cin(gnd),
	.combout(\Mux38~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~17 .lut_mask = 16'hDC98;
defparam \Mux38~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N30
cycloneive_lcell_comb \Mux38~18 (
// Equation(s):
// \Mux38~18_combout  = (instruction_D[17] & ((\Mux38~17_combout  & ((\rfile[15][25]~q ))) # (!\Mux38~17_combout  & (\rfile[14][25]~q )))) # (!instruction_D[17] & (((\Mux38~17_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[14][25]~q ),
	.datac(\rfile[15][25]~q ),
	.datad(\Mux38~17_combout ),
	.cin(gnd),
	.combout(\Mux38~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~18 .lut_mask = 16'hF588;
defparam \Mux38~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N22
cycloneive_lcell_comb \rfile[11][25]~feeder (
// Equation(s):
// \rfile[11][25]~feeder_combout  = \wdat_WB[25]~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[11][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][25]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[11][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N23
dffeas \rfile[11][25] (
	.clk(!CLK),
	.d(\rfile[11][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][25] .is_wysiwyg = "true";
defparam \rfile[11][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N13
dffeas \rfile[9][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][25] .is_wysiwyg = "true";
defparam \rfile[9][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N5
dffeas \rfile[10][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][25] .is_wysiwyg = "true";
defparam \rfile[10][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N27
dffeas \rfile[8][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][25] .is_wysiwyg = "true";
defparam \rfile[8][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N26
cycloneive_lcell_comb \Mux38~10 (
// Equation(s):
// \Mux38~10_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & (\rfile[10][25]~q )) # (!instruction_D[17] & ((\rfile[8][25]~q )))))

	.dataa(instruction_D_16),
	.datab(\rfile[10][25]~q ),
	.datac(\rfile[8][25]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux38~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~10 .lut_mask = 16'hEE50;
defparam \Mux38~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N8
cycloneive_lcell_comb \Mux38~11 (
// Equation(s):
// \Mux38~11_combout  = (instruction_D[16] & ((\Mux38~10_combout  & (\rfile[11][25]~q )) # (!\Mux38~10_combout  & ((\rfile[9][25]~q ))))) # (!instruction_D[16] & (((\Mux38~10_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][25]~q ),
	.datac(\rfile[9][25]~q ),
	.datad(\Mux38~10_combout ),
	.cin(gnd),
	.combout(\Mux38~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~11 .lut_mask = 16'hDDA0;
defparam \Mux38~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N15
dffeas \rfile[7][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][25] .is_wysiwyg = "true";
defparam \rfile[7][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y36_N1
dffeas \rfile[6][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][25] .is_wysiwyg = "true";
defparam \rfile[6][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N5
dffeas \rfile[5][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][25] .is_wysiwyg = "true";
defparam \rfile[5][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N3
dffeas \rfile[4][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][25] .is_wysiwyg = "true";
defparam \rfile[4][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N4
cycloneive_lcell_comb \Mux38~12 (
// Equation(s):
// \Mux38~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[5][25]~q )) # (!instruction_D[16] & ((\rfile[4][25]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[5][25]~q ),
	.datad(\rfile[4][25]~q ),
	.cin(gnd),
	.combout(\Mux38~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~12 .lut_mask = 16'hD9C8;
defparam \Mux38~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N0
cycloneive_lcell_comb \Mux38~13 (
// Equation(s):
// \Mux38~13_combout  = (instruction_D[17] & ((\Mux38~12_combout  & (\rfile[7][25]~q )) # (!\Mux38~12_combout  & ((\rfile[6][25]~q ))))) # (!instruction_D[17] & (((\Mux38~12_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[7][25]~q ),
	.datac(\rfile[6][25]~q ),
	.datad(\Mux38~12_combout ),
	.cin(gnd),
	.combout(\Mux38~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~13 .lut_mask = 16'hDDA0;
defparam \Mux38~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N19
dffeas \rfile[3][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][25] .is_wysiwyg = "true";
defparam \rfile[3][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N29
dffeas \rfile[1][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][25] .is_wysiwyg = "true";
defparam \rfile[1][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N28
cycloneive_lcell_comb \Mux38~14 (
// Equation(s):
// \Mux38~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][25]~q )) # (!instruction_D[17] & ((\rfile[1][25]~q )))))

	.dataa(instruction_D_16),
	.datab(\rfile[3][25]~q ),
	.datac(\rfile[1][25]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux38~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~14 .lut_mask = 16'h88A0;
defparam \Mux38~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N10
cycloneive_lcell_comb \rfile[2][25]~feeder (
// Equation(s):
// \rfile[2][25]~feeder_combout  = \wdat_WB[25]~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_25),
	.cin(gnd),
	.combout(\rfile[2][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][25]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N11
dffeas \rfile[2][25] (
	.clk(!CLK),
	.d(\rfile[2][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][25] .is_wysiwyg = "true";
defparam \rfile[2][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N14
cycloneive_lcell_comb \Mux38~15 (
// Equation(s):
// \Mux38~15_combout  = (\Mux38~14_combout ) # ((instruction_D[17] & (\rfile[2][25]~q  & !instruction_D[16])))

	.dataa(instruction_D_17),
	.datab(\Mux38~14_combout ),
	.datac(\rfile[2][25]~q ),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux38~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~15 .lut_mask = 16'hCCEC;
defparam \Mux38~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N0
cycloneive_lcell_comb \Mux38~16 (
// Equation(s):
// \Mux38~16_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\Mux38~13_combout )))) # (!instruction_D[18] & (!instruction_D[19] & ((\Mux38~15_combout ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\Mux38~13_combout ),
	.datad(\Mux38~15_combout ),
	.cin(gnd),
	.combout(\Mux38~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~16 .lut_mask = 16'hB9A8;
defparam \Mux38~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N15
dffeas \rfile[29][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][24] .is_wysiwyg = "true";
defparam \rfile[29][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N21
dffeas \rfile[21][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][24] .is_wysiwyg = "true";
defparam \rfile[21][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N15
dffeas \rfile[25][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][24] .is_wysiwyg = "true";
defparam \rfile[25][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N25
dffeas \rfile[17][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][24] .is_wysiwyg = "true";
defparam \rfile[17][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N24
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (instruction_D[19] & ((\rfile[25][24]~q ) # ((instruction_D[18])))) # (!instruction_D[19] & (((\rfile[17][24]~q  & !instruction_D[18]))))

	.dataa(instruction_D_19),
	.datab(\rfile[25][24]~q ),
	.datac(\rfile[17][24]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hAAD8;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N20
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (instruction_D[18] & ((\Mux39~0_combout  & (\rfile[29][24]~q )) # (!\Mux39~0_combout  & ((\rfile[21][24]~q ))))) # (!instruction_D[18] & (((\Mux39~0_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[29][24]~q ),
	.datac(\rfile[21][24]~q ),
	.datad(\Mux39~0_combout ),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hDDA0;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y35_N17
dffeas \rfile[18][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][24] .is_wysiwyg = "true";
defparam \rfile[18][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y35_N31
dffeas \rfile[22][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][24] .is_wysiwyg = "true";
defparam \rfile[22][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N16
cycloneive_lcell_comb \Mux39~2 (
// Equation(s):
// \Mux39~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[22][24]~q ))) # (!instruction_D[18] & (\rfile[18][24]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][24]~q ),
	.datad(\rfile[22][24]~q ),
	.cin(gnd),
	.combout(\Mux39~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~2 .lut_mask = 16'hDC98;
defparam \Mux39~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y34_N1
dffeas \rfile[30][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][24] .is_wysiwyg = "true";
defparam \rfile[30][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y34_N19
dffeas \rfile[26][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][24] .is_wysiwyg = "true";
defparam \rfile[26][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N0
cycloneive_lcell_comb \Mux39~3 (
// Equation(s):
// \Mux39~3_combout  = (instruction_D[19] & ((\Mux39~2_combout  & (\rfile[30][24]~q )) # (!\Mux39~2_combout  & ((\rfile[26][24]~q ))))) # (!instruction_D[19] & (\Mux39~2_combout ))

	.dataa(instruction_D_19),
	.datab(\Mux39~2_combout ),
	.datac(\rfile[30][24]~q ),
	.datad(\rfile[26][24]~q ),
	.cin(gnd),
	.combout(\Mux39~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~3 .lut_mask = 16'hE6C4;
defparam \Mux39~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N31
dffeas \rfile[28][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][24] .is_wysiwyg = "true";
defparam \rfile[28][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N29
dffeas \rfile[24][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][24] .is_wysiwyg = "true";
defparam \rfile[24][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N30
cycloneive_lcell_comb \Mux39~5 (
// Equation(s):
// \Mux39~5_combout  = (\Mux39~4_combout  & (((\rfile[28][24]~q )) # (!instruction_D[19]))) # (!\Mux39~4_combout  & (instruction_D[19] & ((\rfile[24][24]~q ))))

	.dataa(\Mux39~4_combout ),
	.datab(instruction_D_19),
	.datac(\rfile[28][24]~q ),
	.datad(\rfile[24][24]~q ),
	.cin(gnd),
	.combout(\Mux39~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~5 .lut_mask = 16'hE6A2;
defparam \Mux39~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N4
cycloneive_lcell_comb \Mux39~6 (
// Equation(s):
// \Mux39~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\Mux39~3_combout )) # (!instruction_D[17] & ((\Mux39~5_combout )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux39~3_combout ),
	.datad(\Mux39~5_combout ),
	.cin(gnd),
	.combout(\Mux39~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~6 .lut_mask = 16'hD9C8;
defparam \Mux39~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N8
cycloneive_lcell_comb \rfile[23][24]~feeder (
// Equation(s):
// \rfile[23][24]~feeder_combout  = \wdat_WB[24]~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_24),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[23][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[23][24]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[23][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N9
dffeas \rfile[23][24] (
	.clk(!CLK),
	.d(\rfile[23][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][24] .is_wysiwyg = "true";
defparam \rfile[23][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N7
dffeas \rfile[31][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][24] .is_wysiwyg = "true";
defparam \rfile[31][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N5
dffeas \rfile[27][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][24] .is_wysiwyg = "true";
defparam \rfile[27][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N23
dffeas \rfile[19][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][24] .is_wysiwyg = "true";
defparam \rfile[19][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N22
cycloneive_lcell_comb \Mux39~7 (
// Equation(s):
// \Mux39~7_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[27][24]~q )) # (!instruction_D[19] & ((\rfile[19][24]~q )))))

	.dataa(instruction_D_18),
	.datab(\rfile[27][24]~q ),
	.datac(\rfile[19][24]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux39~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~7 .lut_mask = 16'hEE50;
defparam \Mux39~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N6
cycloneive_lcell_comb \Mux39~8 (
// Equation(s):
// \Mux39~8_combout  = (instruction_D[18] & ((\Mux39~7_combout  & ((\rfile[31][24]~q ))) # (!\Mux39~7_combout  & (\rfile[23][24]~q )))) # (!instruction_D[18] & (((\Mux39~7_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[23][24]~q ),
	.datac(\rfile[31][24]~q ),
	.datad(\Mux39~7_combout ),
	.cin(gnd),
	.combout(\Mux39~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~8 .lut_mask = 16'hF588;
defparam \Mux39~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N23
dffeas \rfile[7][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][24] .is_wysiwyg = "true";
defparam \rfile[7][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N4
cycloneive_lcell_comb \rfile[6][24]~feeder (
// Equation(s):
// \rfile[6][24]~feeder_combout  = \wdat_WB[24]~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_24),
	.cin(gnd),
	.combout(\rfile[6][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][24]~feeder .lut_mask = 16'hFF00;
defparam \rfile[6][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N5
dffeas \rfile[6][24] (
	.clk(!CLK),
	.d(\rfile[6][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][24] .is_wysiwyg = "true";
defparam \rfile[6][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N1
dffeas \rfile[5][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][24] .is_wysiwyg = "true";
defparam \rfile[5][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N0
cycloneive_lcell_comb \Mux39~10 (
// Equation(s):
// \Mux39~10_combout  = (instruction_D[16] & (((\rfile[5][24]~q ) # (instruction_D[17])))) # (!instruction_D[16] & (\rfile[4][24]~q  & ((!instruction_D[17]))))

	.dataa(\rfile[4][24]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[5][24]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux39~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~10 .lut_mask = 16'hCCE2;
defparam \Mux39~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N16
cycloneive_lcell_comb \Mux39~11 (
// Equation(s):
// \Mux39~11_combout  = (instruction_D[17] & ((\Mux39~10_combout  & (\rfile[7][24]~q )) # (!\Mux39~10_combout  & ((\rfile[6][24]~q ))))) # (!instruction_D[17] & (((\Mux39~10_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[7][24]~q ),
	.datac(\rfile[6][24]~q ),
	.datad(\Mux39~10_combout ),
	.cin(gnd),
	.combout(\Mux39~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~11 .lut_mask = 16'hDDA0;
defparam \Mux39~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N20
cycloneive_lcell_comb \rfile[2][24]~feeder (
// Equation(s):
// \rfile[2][24]~feeder_combout  = \wdat_WB[24]~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_24),
	.cin(gnd),
	.combout(\rfile[2][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][24]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N21
dffeas \rfile[2][24] (
	.clk(!CLK),
	.d(\rfile[2][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][24] .is_wysiwyg = "true";
defparam \rfile[2][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N11
dffeas \rfile[1][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][24] .is_wysiwyg = "true";
defparam \rfile[1][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N21
dffeas \rfile[3][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][24] .is_wysiwyg = "true";
defparam \rfile[3][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N10
cycloneive_lcell_comb \Mux39~14 (
// Equation(s):
// \Mux39~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][24]~q ))) # (!instruction_D[17] & (\rfile[1][24]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[1][24]~q ),
	.datad(\rfile[3][24]~q ),
	.cin(gnd),
	.combout(\Mux39~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~14 .lut_mask = 16'hC840;
defparam \Mux39~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N4
cycloneive_lcell_comb \Mux39~15 (
// Equation(s):
// \Mux39~15_combout  = (\Mux39~14_combout ) # ((!instruction_D[16] & (\rfile[2][24]~q  & instruction_D[17])))

	.dataa(instruction_D_16),
	.datab(\rfile[2][24]~q ),
	.datac(\Mux39~14_combout ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux39~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~15 .lut_mask = 16'hF4F0;
defparam \Mux39~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N0
cycloneive_lcell_comb \rfile[11][24]~feeder (
// Equation(s):
// \rfile[11][24]~feeder_combout  = \wdat_WB[24]~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_24),
	.cin(gnd),
	.combout(\rfile[11][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][24]~feeder .lut_mask = 16'hFF00;
defparam \rfile[11][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N1
dffeas \rfile[11][24] (
	.clk(!CLK),
	.d(\rfile[11][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][24] .is_wysiwyg = "true";
defparam \rfile[11][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N23
dffeas \rfile[8][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][24] .is_wysiwyg = "true";
defparam \rfile[8][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N1
dffeas \rfile[10][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][24] .is_wysiwyg = "true";
defparam \rfile[10][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N22
cycloneive_lcell_comb \Mux39~12 (
// Equation(s):
// \Mux39~12_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][24]~q ))) # (!instruction_D[17] & (\rfile[8][24]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[8][24]~q ),
	.datad(\rfile[10][24]~q ),
	.cin(gnd),
	.combout(\Mux39~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~12 .lut_mask = 16'hDC98;
defparam \Mux39~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N14
cycloneive_lcell_comb \Mux39~13 (
// Equation(s):
// \Mux39~13_combout  = (instruction_D[16] & ((\Mux39~12_combout  & ((\rfile[11][24]~q ))) # (!\Mux39~12_combout  & (\rfile[9][24]~q )))) # (!instruction_D[16] & (((\Mux39~12_combout ))))

	.dataa(\rfile[9][24]~q ),
	.datab(\rfile[11][24]~q ),
	.datac(instruction_D_16),
	.datad(\Mux39~12_combout ),
	.cin(gnd),
	.combout(\Mux39~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~13 .lut_mask = 16'hCFA0;
defparam \Mux39~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N14
cycloneive_lcell_comb \Mux39~16 (
// Equation(s):
// \Mux39~16_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\Mux39~13_combout ))) # (!instruction_D[19] & (\Mux39~15_combout ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\Mux39~15_combout ),
	.datad(\Mux39~13_combout ),
	.cin(gnd),
	.combout(\Mux39~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~16 .lut_mask = 16'hDC98;
defparam \Mux39~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N20
cycloneive_lcell_comb \rfile[15][24]~feeder (
// Equation(s):
// \rfile[15][24]~feeder_combout  = \wdat_WB[24]~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_24),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[15][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][24]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[15][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N21
dffeas \rfile[15][24] (
	.clk(!CLK),
	.d(\rfile[15][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][24] .is_wysiwyg = "true";
defparam \rfile[15][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N19
dffeas \rfile[14][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][24] .is_wysiwyg = "true";
defparam \rfile[14][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N27
dffeas \rfile[12][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][24] .is_wysiwyg = "true";
defparam \rfile[12][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N18
cycloneive_lcell_comb \rfile[13][24]~feeder (
// Equation(s):
// \rfile[13][24]~feeder_combout  = \wdat_WB[24]~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_24),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[13][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[13][24]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[13][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N19
dffeas \rfile[13][24] (
	.clk(!CLK),
	.d(\rfile[13][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][24] .is_wysiwyg = "true";
defparam \rfile[13][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N16
cycloneive_lcell_comb \Mux39~17 (
// Equation(s):
// \Mux39~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][24]~q ))) # (!instruction_D[16] & (\rfile[12][24]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][24]~q ),
	.datad(\rfile[13][24]~q ),
	.cin(gnd),
	.combout(\Mux39~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~17 .lut_mask = 16'hDC98;
defparam \Mux39~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N18
cycloneive_lcell_comb \Mux39~18 (
// Equation(s):
// \Mux39~18_combout  = (instruction_D[17] & ((\Mux39~17_combout  & (\rfile[15][24]~q )) # (!\Mux39~17_combout  & ((\rfile[14][24]~q ))))) # (!instruction_D[17] & (((\Mux39~17_combout ))))

	.dataa(\rfile[15][24]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[14][24]~q ),
	.datad(\Mux39~17_combout ),
	.cin(gnd),
	.combout(\Mux39~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~18 .lut_mask = 16'hBBC0;
defparam \Mux39~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N16
cycloneive_lcell_comb \rfile[25][23]~feeder (
// Equation(s):
// \rfile[25][23]~feeder_combout  = \wdat_WB[23]~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_23),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[25][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[25][23]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[25][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N17
dffeas \rfile[25][23] (
	.clk(!CLK),
	.d(\rfile[25][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][23] .is_wysiwyg = "true";
defparam \rfile[25][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N29
dffeas \rfile[29][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][23] .is_wysiwyg = "true";
defparam \rfile[29][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N5
dffeas \rfile[21][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][23] .is_wysiwyg = "true";
defparam \rfile[21][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N30
cycloneive_lcell_comb \rfile[17][23]~feeder (
// Equation(s):
// \rfile[17][23]~feeder_combout  = \wdat_WB[23]~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_23),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[17][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[17][23]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[17][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y27_N31
dffeas \rfile[17][23] (
	.clk(!CLK),
	.d(\rfile[17][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][23] .is_wysiwyg = "true";
defparam \rfile[17][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N18
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[21][23]~q )) # (!instruction_D[18] & ((\rfile[17][23]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[21][23]~q ),
	.datad(\rfile[17][23]~q ),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hD9C8;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N28
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (instruction_D[19] & ((\Mux40~0_combout  & ((\rfile[29][23]~q ))) # (!\Mux40~0_combout  & (\rfile[25][23]~q )))) # (!instruction_D[19] & (((\Mux40~0_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[25][23]~q ),
	.datac(\rfile[29][23]~q ),
	.datad(\Mux40~0_combout ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hF588;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y28_N29
dffeas \rfile[27][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][23] .is_wysiwyg = "true";
defparam \rfile[27][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N19
dffeas \rfile[31][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][23] .is_wysiwyg = "true";
defparam \rfile[31][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N27
dffeas \rfile[19][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][23] .is_wysiwyg = "true";
defparam \rfile[19][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N13
dffeas \rfile[23][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][23] .is_wysiwyg = "true";
defparam \rfile[23][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N26
cycloneive_lcell_comb \Mux40~7 (
// Equation(s):
// \Mux40~7_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[23][23]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[19][23]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[19][23]~q ),
	.datad(\rfile[23][23]~q ),
	.cin(gnd),
	.combout(\Mux40~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~7 .lut_mask = 16'hBA98;
defparam \Mux40~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N18
cycloneive_lcell_comb \Mux40~8 (
// Equation(s):
// \Mux40~8_combout  = (instruction_D[19] & ((\Mux40~7_combout  & ((\rfile[31][23]~q ))) # (!\Mux40~7_combout  & (\rfile[27][23]~q )))) # (!instruction_D[19] & (((\Mux40~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[27][23]~q ),
	.datac(\rfile[31][23]~q ),
	.datad(\Mux40~7_combout ),
	.cin(gnd),
	.combout(\Mux40~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~8 .lut_mask = 16'hF588;
defparam \Mux40~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N8
cycloneive_lcell_comb \rfile[20][23]~feeder (
// Equation(s):
// \rfile[20][23]~feeder_combout  = \wdat_WB[23]~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_23),
	.cin(gnd),
	.combout(\rfile[20][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[20][23]~feeder .lut_mask = 16'hFF00;
defparam \rfile[20][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y31_N9
dffeas \rfile[20][23] (
	.clk(!CLK),
	.d(\rfile[20][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][23] .is_wysiwyg = "true";
defparam \rfile[20][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N5
dffeas \rfile[28][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][23] .is_wysiwyg = "true";
defparam \rfile[28][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y32_N25
dffeas \rfile[16][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][23] .is_wysiwyg = "true";
defparam \rfile[16][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y32_N13
dffeas \rfile[24][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][23] .is_wysiwyg = "true";
defparam \rfile[24][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N24
cycloneive_lcell_comb \Mux40~4 (
// Equation(s):
// \Mux40~4_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[24][23]~q )))) # (!instruction_D[19] & (!instruction_D[18] & (\rfile[16][23]~q )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[16][23]~q ),
	.datad(\rfile[24][23]~q ),
	.cin(gnd),
	.combout(\Mux40~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~4 .lut_mask = 16'hBA98;
defparam \Mux40~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N4
cycloneive_lcell_comb \Mux40~5 (
// Equation(s):
// \Mux40~5_combout  = (instruction_D[18] & ((\Mux40~4_combout  & ((\rfile[28][23]~q ))) # (!\Mux40~4_combout  & (\rfile[20][23]~q )))) # (!instruction_D[18] & (((\Mux40~4_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[20][23]~q ),
	.datac(\rfile[28][23]~q ),
	.datad(\Mux40~4_combout ),
	.cin(gnd),
	.combout(\Mux40~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~5 .lut_mask = 16'hF588;
defparam \Mux40~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N0
cycloneive_lcell_comb \rfile[22][23]~feeder (
// Equation(s):
// \rfile[22][23]~feeder_combout  = \wdat_WB[23]~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_23),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[22][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[22][23]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[22][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N1
dffeas \rfile[22][23] (
	.clk(!CLK),
	.d(\rfile[22][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][23] .is_wysiwyg = "true";
defparam \rfile[22][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y34_N31
dffeas \rfile[30][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][23] .is_wysiwyg = "true";
defparam \rfile[30][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y34_N25
dffeas \rfile[18][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][23] .is_wysiwyg = "true";
defparam \rfile[18][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N18
cycloneive_lcell_comb \rfile[26][23]~feeder (
// Equation(s):
// \rfile[26][23]~feeder_combout  = \wdat_WB[23]~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_23),
	.cin(gnd),
	.combout(\rfile[26][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[26][23]~feeder .lut_mask = 16'hFF00;
defparam \rfile[26][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y36_N19
dffeas \rfile[26][23] (
	.clk(!CLK),
	.d(\rfile[26][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][23] .is_wysiwyg = "true";
defparam \rfile[26][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N24
cycloneive_lcell_comb \Mux40~2 (
// Equation(s):
// \Mux40~2_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[26][23]~q )))) # (!instruction_D[19] & (!instruction_D[18] & (\rfile[18][23]~q )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][23]~q ),
	.datad(\rfile[26][23]~q ),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~2 .lut_mask = 16'hBA98;
defparam \Mux40~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N30
cycloneive_lcell_comb \Mux40~3 (
// Equation(s):
// \Mux40~3_combout  = (instruction_D[18] & ((\Mux40~2_combout  & ((\rfile[30][23]~q ))) # (!\Mux40~2_combout  & (\rfile[22][23]~q )))) # (!instruction_D[18] & (((\Mux40~2_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[22][23]~q ),
	.datac(\rfile[30][23]~q ),
	.datad(\Mux40~2_combout ),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~3 .lut_mask = 16'hF588;
defparam \Mux40~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N20
cycloneive_lcell_comb \Mux40~6 (
// Equation(s):
// \Mux40~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\Mux40~3_combout ))) # (!instruction_D[17] & (\Mux40~5_combout ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux40~5_combout ),
	.datad(\Mux40~3_combout ),
	.cin(gnd),
	.combout(\Mux40~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~6 .lut_mask = 16'hDC98;
defparam \Mux40~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N0
cycloneive_lcell_comb \rfile[2][23]~feeder (
// Equation(s):
// \rfile[2][23]~feeder_combout  = \wdat_WB[23]~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_23),
	.cin(gnd),
	.combout(\rfile[2][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][23]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N1
dffeas \rfile[2][23] (
	.clk(!CLK),
	.d(\rfile[2][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][23] .is_wysiwyg = "true";
defparam \rfile[2][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N25
dffeas \rfile[3][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][23] .is_wysiwyg = "true";
defparam \rfile[3][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N19
dffeas \rfile[1][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][23] .is_wysiwyg = "true";
defparam \rfile[1][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N24
cycloneive_lcell_comb \Mux40~14 (
// Equation(s):
// \Mux40~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][23]~q )) # (!instruction_D[17] & ((\rfile[1][23]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[3][23]~q ),
	.datad(\rfile[1][23]~q ),
	.cin(gnd),
	.combout(\Mux40~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~14 .lut_mask = 16'hC480;
defparam \Mux40~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N26
cycloneive_lcell_comb \Mux40~15 (
// Equation(s):
// \Mux40~15_combout  = (\Mux40~14_combout ) # ((!instruction_D[16] & (\rfile[2][23]~q  & instruction_D[17])))

	.dataa(instruction_D_16),
	.datab(\rfile[2][23]~q ),
	.datac(instruction_D_17),
	.datad(\Mux40~14_combout ),
	.cin(gnd),
	.combout(\Mux40~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~15 .lut_mask = 16'hFF40;
defparam \Mux40~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N3
dffeas \rfile[7][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][23] .is_wysiwyg = "true";
defparam \rfile[7][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N15
dffeas \rfile[5][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][23] .is_wysiwyg = "true";
defparam \rfile[5][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y28_N25
dffeas \rfile[4][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][23] .is_wysiwyg = "true";
defparam \rfile[4][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N14
cycloneive_lcell_comb \Mux40~12 (
// Equation(s):
// \Mux40~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[5][23]~q )) # (!instruction_D[16] & ((\rfile[4][23]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[5][23]~q ),
	.datad(\rfile[4][23]~q ),
	.cin(gnd),
	.combout(\Mux40~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~12 .lut_mask = 16'hD9C8;
defparam \Mux40~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N10
cycloneive_lcell_comb \Mux40~13 (
// Equation(s):
// \Mux40~13_combout  = (instruction_D[17] & ((\Mux40~12_combout  & ((\rfile[7][23]~q ))) # (!\Mux40~12_combout  & (\rfile[6][23]~q )))) # (!instruction_D[17] & (((\Mux40~12_combout ))))

	.dataa(\rfile[6][23]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[7][23]~q ),
	.datad(\Mux40~12_combout ),
	.cin(gnd),
	.combout(\Mux40~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~13 .lut_mask = 16'hF388;
defparam \Mux40~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N24
cycloneive_lcell_comb \Mux40~16 (
// Equation(s):
// \Mux40~16_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\Mux40~13_combout ))) # (!instruction_D[18] & (\Mux40~15_combout ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux40~15_combout ),
	.datad(\Mux40~13_combout ),
	.cin(gnd),
	.combout(\Mux40~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~16 .lut_mask = 16'hDC98;
defparam \Mux40~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N23
dffeas \rfile[11][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][23] .is_wysiwyg = "true";
defparam \rfile[11][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N1
dffeas \rfile[9][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][23] .is_wysiwyg = "true";
defparam \rfile[9][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N31
dffeas \rfile[8][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][23] .is_wysiwyg = "true";
defparam \rfile[8][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N25
dffeas \rfile[10][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][23] .is_wysiwyg = "true";
defparam \rfile[10][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N30
cycloneive_lcell_comb \Mux40~10 (
// Equation(s):
// \Mux40~10_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][23]~q )))) # (!instruction_D[17] & (!instruction_D[16] & (\rfile[8][23]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[8][23]~q ),
	.datad(\rfile[10][23]~q ),
	.cin(gnd),
	.combout(\Mux40~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~10 .lut_mask = 16'hBA98;
defparam \Mux40~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N0
cycloneive_lcell_comb \Mux40~11 (
// Equation(s):
// \Mux40~11_combout  = (instruction_D[16] & ((\Mux40~10_combout  & (\rfile[11][23]~q )) # (!\Mux40~10_combout  & ((\rfile[9][23]~q ))))) # (!instruction_D[16] & (((\Mux40~10_combout ))))

	.dataa(\rfile[11][23]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[9][23]~q ),
	.datad(\Mux40~10_combout ),
	.cin(gnd),
	.combout(\Mux40~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~11 .lut_mask = 16'hBBC0;
defparam \Mux40~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N5
dffeas \rfile[13][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][23] .is_wysiwyg = "true";
defparam \rfile[13][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N3
dffeas \rfile[12][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][23] .is_wysiwyg = "true";
defparam \rfile[12][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N4
cycloneive_lcell_comb \Mux40~17 (
// Equation(s):
// \Mux40~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[13][23]~q )) # (!instruction_D[16] & ((\rfile[12][23]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[13][23]~q ),
	.datad(\rfile[12][23]~q ),
	.cin(gnd),
	.combout(\Mux40~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~17 .lut_mask = 16'hD9C8;
defparam \Mux40~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N3
dffeas \rfile[14][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][23] .is_wysiwyg = "true";
defparam \rfile[14][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N20
cycloneive_lcell_comb \rfile[15][23]~feeder (
// Equation(s):
// \rfile[15][23]~feeder_combout  = \wdat_WB[23]~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_23),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[15][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][23]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[15][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N21
dffeas \rfile[15][23] (
	.clk(!CLK),
	.d(\rfile[15][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][23] .is_wysiwyg = "true";
defparam \rfile[15][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N2
cycloneive_lcell_comb \Mux40~18 (
// Equation(s):
// \Mux40~18_combout  = (\Mux40~17_combout  & (((\rfile[15][23]~q )) # (!instruction_D[17]))) # (!\Mux40~17_combout  & (instruction_D[17] & (\rfile[14][23]~q )))

	.dataa(\Mux40~17_combout ),
	.datab(instruction_D_17),
	.datac(\rfile[14][23]~q ),
	.datad(\rfile[15][23]~q ),
	.cin(gnd),
	.combout(\Mux40~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~18 .lut_mask = 16'hEA62;
defparam \Mux40~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N12
cycloneive_lcell_comb \rfile[29][22]~feeder (
// Equation(s):
// \rfile[29][22]~feeder_combout  = \wdat_WB[22]~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[29][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[29][22]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[29][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N13
dffeas \rfile[29][22] (
	.clk(!CLK),
	.d(\rfile[29][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][22] .is_wysiwyg = "true";
defparam \rfile[29][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N31
dffeas \rfile[21][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][22] .is_wysiwyg = "true";
defparam \rfile[21][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N11
dffeas \rfile[17][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][22] .is_wysiwyg = "true";
defparam \rfile[17][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N13
dffeas \rfile[25][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][22] .is_wysiwyg = "true";
defparam \rfile[25][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N10
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[25][22]~q )))) # (!instruction_D[19] & (!instruction_D[18] & (\rfile[17][22]~q )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[17][22]~q ),
	.datad(\rfile[25][22]~q ),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hBA98;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N30
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (instruction_D[18] & ((\Mux41~0_combout  & (\rfile[29][22]~q )) # (!\Mux41~0_combout  & ((\rfile[21][22]~q ))))) # (!instruction_D[18] & (((\Mux41~0_combout ))))

	.dataa(\rfile[29][22]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[21][22]~q ),
	.datad(\Mux41~0_combout ),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hBBC0;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y28_N19
dffeas \rfile[19][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][22] .is_wysiwyg = "true";
defparam \rfile[19][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N13
dffeas \rfile[27][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][22] .is_wysiwyg = "true";
defparam \rfile[27][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N18
cycloneive_lcell_comb \Mux41~7 (
// Equation(s):
// \Mux41~7_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[27][22]~q ))) # (!instruction_D[19] & (\rfile[19][22]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[19][22]~q ),
	.datad(\rfile[27][22]~q ),
	.cin(gnd),
	.combout(\Mux41~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~7 .lut_mask = 16'hDC98;
defparam \Mux41~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N15
dffeas \rfile[31][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][22] .is_wysiwyg = "true";
defparam \rfile[31][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N1
dffeas \rfile[23][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][22] .is_wysiwyg = "true";
defparam \rfile[23][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N14
cycloneive_lcell_comb \Mux41~8 (
// Equation(s):
// \Mux41~8_combout  = (instruction_D[18] & ((\Mux41~7_combout  & (\rfile[31][22]~q )) # (!\Mux41~7_combout  & ((\rfile[23][22]~q ))))) # (!instruction_D[18] & (\Mux41~7_combout ))

	.dataa(instruction_D_18),
	.datab(\Mux41~7_combout ),
	.datac(\rfile[31][22]~q ),
	.datad(\rfile[23][22]~q ),
	.cin(gnd),
	.combout(\Mux41~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~8 .lut_mask = 16'hE6C4;
defparam \Mux41~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N8
cycloneive_lcell_comb \rfile[24][22]~feeder (
// Equation(s):
// \rfile[24][22]~feeder_combout  = \wdat_WB[22]~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[24][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[24][22]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[24][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y30_N9
dffeas \rfile[24][22] (
	.clk(!CLK),
	.d(\rfile[24][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][22] .is_wysiwyg = "true";
defparam \rfile[24][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y31_N25
dffeas \rfile[16][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][22] .is_wysiwyg = "true";
defparam \rfile[16][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y31_N7
dffeas \rfile[20][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][22] .is_wysiwyg = "true";
defparam \rfile[20][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N24
cycloneive_lcell_comb \Mux41~4 (
// Equation(s):
// \Mux41~4_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[20][22]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[16][22]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[16][22]~q ),
	.datad(\rfile[20][22]~q ),
	.cin(gnd),
	.combout(\Mux41~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~4 .lut_mask = 16'hBA98;
defparam \Mux41~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N0
cycloneive_lcell_comb \Mux41~5 (
// Equation(s):
// \Mux41~5_combout  = (instruction_D[19] & ((\Mux41~4_combout  & (\rfile[28][22]~q )) # (!\Mux41~4_combout  & ((\rfile[24][22]~q ))))) # (!instruction_D[19] & (((\Mux41~4_combout ))))

	.dataa(\rfile[28][22]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[24][22]~q ),
	.datad(\Mux41~4_combout ),
	.cin(gnd),
	.combout(\Mux41~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~5 .lut_mask = 16'hBBC0;
defparam \Mux41~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y34_N25
dffeas \rfile[30][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][22] .is_wysiwyg = "true";
defparam \rfile[30][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y34_N27
dffeas \rfile[26][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][22] .is_wysiwyg = "true";
defparam \rfile[26][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y34_N27
dffeas \rfile[22][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][22] .is_wysiwyg = "true";
defparam \rfile[22][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y34_N29
dffeas \rfile[18][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][22] .is_wysiwyg = "true";
defparam \rfile[18][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N26
cycloneive_lcell_comb \Mux41~2 (
// Equation(s):
// \Mux41~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[22][22]~q )) # (!instruction_D[18] & ((\rfile[18][22]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[22][22]~q ),
	.datad(\rfile[18][22]~q ),
	.cin(gnd),
	.combout(\Mux41~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~2 .lut_mask = 16'hD9C8;
defparam \Mux41~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N26
cycloneive_lcell_comb \Mux41~3 (
// Equation(s):
// \Mux41~3_combout  = (instruction_D[19] & ((\Mux41~2_combout  & (\rfile[30][22]~q )) # (!\Mux41~2_combout  & ((\rfile[26][22]~q ))))) # (!instruction_D[19] & (((\Mux41~2_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[30][22]~q ),
	.datac(\rfile[26][22]~q ),
	.datad(\Mux41~2_combout ),
	.cin(gnd),
	.combout(\Mux41~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~3 .lut_mask = 16'hDDA0;
defparam \Mux41~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N0
cycloneive_lcell_comb \Mux41~6 (
// Equation(s):
// \Mux41~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux41~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & (\Mux41~5_combout )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux41~5_combout ),
	.datad(\Mux41~3_combout ),
	.cin(gnd),
	.combout(\Mux41~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~6 .lut_mask = 16'hBA98;
defparam \Mux41~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N24
cycloneive_lcell_comb \rfile[14][22]~feeder (
// Equation(s):
// \rfile[14][22]~feeder_combout  = \wdat_WB[22]~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[14][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][22]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[14][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N25
dffeas \rfile[14][22] (
	.clk(!CLK),
	.d(\rfile[14][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][22] .is_wysiwyg = "true";
defparam \rfile[14][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N21
dffeas \rfile[13][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][22] .is_wysiwyg = "true";
defparam \rfile[13][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N19
dffeas \rfile[12][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][22] .is_wysiwyg = "true";
defparam \rfile[12][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N20
cycloneive_lcell_comb \Mux41~17 (
// Equation(s):
// \Mux41~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[13][22]~q )) # (!instruction_D[16] & ((\rfile[12][22]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[13][22]~q ),
	.datad(\rfile[12][22]~q ),
	.cin(gnd),
	.combout(\Mux41~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~17 .lut_mask = 16'hD9C8;
defparam \Mux41~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N26
cycloneive_lcell_comb \rfile[15][22]~feeder (
// Equation(s):
// \rfile[15][22]~feeder_combout  = \wdat_WB[22]~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[15][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][22]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[15][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N27
dffeas \rfile[15][22] (
	.clk(!CLK),
	.d(\rfile[15][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][22] .is_wysiwyg = "true";
defparam \rfile[15][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N26
cycloneive_lcell_comb \Mux41~18 (
// Equation(s):
// \Mux41~18_combout  = (instruction_D[17] & ((\Mux41~17_combout  & ((\rfile[15][22]~q ))) # (!\Mux41~17_combout  & (\rfile[14][22]~q )))) # (!instruction_D[17] & (((\Mux41~17_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[14][22]~q ),
	.datac(\Mux41~17_combout ),
	.datad(\rfile[15][22]~q ),
	.cin(gnd),
	.combout(\Mux41~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~18 .lut_mask = 16'hF858;
defparam \Mux41~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N9
dffeas \rfile[2][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][22] .is_wysiwyg = "true";
defparam \rfile[2][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N29
dffeas \rfile[1][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][22] .is_wysiwyg = "true";
defparam \rfile[1][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N3
dffeas \rfile[3][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][22] .is_wysiwyg = "true";
defparam \rfile[3][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N28
cycloneive_lcell_comb \Mux41~14 (
// Equation(s):
// \Mux41~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][22]~q ))) # (!instruction_D[17] & (\rfile[1][22]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[1][22]~q ),
	.datad(\rfile[3][22]~q ),
	.cin(gnd),
	.combout(\Mux41~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~14 .lut_mask = 16'hC840;
defparam \Mux41~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N22
cycloneive_lcell_comb \Mux41~15 (
// Equation(s):
// \Mux41~15_combout  = (\Mux41~14_combout ) # ((instruction_D[17] & (!instruction_D[16] & \rfile[2][22]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[2][22]~q ),
	.datad(\Mux41~14_combout ),
	.cin(gnd),
	.combout(\Mux41~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~15 .lut_mask = 16'hFF20;
defparam \Mux41~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N16
cycloneive_lcell_comb \rfile[11][22]~feeder (
// Equation(s):
// \rfile[11][22]~feeder_combout  = \wdat_WB[22]~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_22),
	.cin(gnd),
	.combout(\rfile[11][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][22]~feeder .lut_mask = 16'hFF00;
defparam \rfile[11][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N17
dffeas \rfile[11][22] (
	.clk(!CLK),
	.d(\rfile[11][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][22] .is_wysiwyg = "true";
defparam \rfile[11][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y35_N27
dffeas \rfile[9][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][22] .is_wysiwyg = "true";
defparam \rfile[9][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N11
dffeas \rfile[8][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][22] .is_wysiwyg = "true";
defparam \rfile[8][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N29
dffeas \rfile[10][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][22] .is_wysiwyg = "true";
defparam \rfile[10][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N10
cycloneive_lcell_comb \Mux41~12 (
// Equation(s):
// \Mux41~12_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][22]~q )))) # (!instruction_D[17] & (!instruction_D[16] & (\rfile[8][22]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[8][22]~q ),
	.datad(\rfile[10][22]~q ),
	.cin(gnd),
	.combout(\Mux41~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~12 .lut_mask = 16'hBA98;
defparam \Mux41~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N26
cycloneive_lcell_comb \Mux41~13 (
// Equation(s):
// \Mux41~13_combout  = (instruction_D[16] & ((\Mux41~12_combout  & (\rfile[11][22]~q )) # (!\Mux41~12_combout  & ((\rfile[9][22]~q ))))) # (!instruction_D[16] & (((\Mux41~12_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][22]~q ),
	.datac(\rfile[9][22]~q ),
	.datad(\Mux41~12_combout ),
	.cin(gnd),
	.combout(\Mux41~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~13 .lut_mask = 16'hDDA0;
defparam \Mux41~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N8
cycloneive_lcell_comb \Mux41~16 (
// Equation(s):
// \Mux41~16_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\Mux41~13_combout )))) # (!instruction_D[19] & (!instruction_D[18] & (\Mux41~15_combout )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux41~15_combout ),
	.datad(\Mux41~13_combout ),
	.cin(gnd),
	.combout(\Mux41~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~16 .lut_mask = 16'hBA98;
defparam \Mux41~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N12
cycloneive_lcell_comb \rfile[6][22]~feeder (
// Equation(s):
// \rfile[6][22]~feeder_combout  = \wdat_WB[22]~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_22),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[6][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][22]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[6][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y27_N13
dffeas \rfile[6][22] (
	.clk(!CLK),
	.d(\rfile[6][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][22] .is_wysiwyg = "true";
defparam \rfile[6][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N11
dffeas \rfile[7][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][22] .is_wysiwyg = "true";
defparam \rfile[7][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N7
dffeas \rfile[4][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][22] .is_wysiwyg = "true";
defparam \rfile[4][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N25
dffeas \rfile[5][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][22] .is_wysiwyg = "true";
defparam \rfile[5][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N6
cycloneive_lcell_comb \Mux41~10 (
// Equation(s):
// \Mux41~10_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][22]~q ))) # (!instruction_D[16] & (\rfile[4][22]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][22]~q ),
	.datad(\rfile[5][22]~q ),
	.cin(gnd),
	.combout(\Mux41~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~10 .lut_mask = 16'hDC98;
defparam \Mux41~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N12
cycloneive_lcell_comb \Mux41~11 (
// Equation(s):
// \Mux41~11_combout  = (instruction_D[17] & ((\Mux41~10_combout  & ((\rfile[7][22]~q ))) # (!\Mux41~10_combout  & (\rfile[6][22]~q )))) # (!instruction_D[17] & (((\Mux41~10_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[6][22]~q ),
	.datac(\rfile[7][22]~q ),
	.datad(\Mux41~10_combout ),
	.cin(gnd),
	.combout(\Mux41~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~11 .lut_mask = 16'hF588;
defparam \Mux41~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N9
dffeas \rfile[29][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][21] .is_wysiwyg = "true";
defparam \rfile[29][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N19
dffeas \rfile[25][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][21] .is_wysiwyg = "true";
defparam \rfile[25][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N17
dffeas \rfile[21][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][21] .is_wysiwyg = "true";
defparam \rfile[21][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N29
dffeas \rfile[17][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][21] .is_wysiwyg = "true";
defparam \rfile[17][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N16
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[21][21]~q )) # (!instruction_D[18] & ((\rfile[17][21]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[21][21]~q ),
	.datad(\rfile[17][21]~q ),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hD9C8;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N18
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (instruction_D[19] & ((\Mux42~0_combout  & (\rfile[29][21]~q )) # (!\Mux42~0_combout  & ((\rfile[25][21]~q ))))) # (!instruction_D[19] & (((\Mux42~0_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[29][21]~q ),
	.datac(\rfile[25][21]~q ),
	.datad(\Mux42~0_combout ),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hDDA0;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y28_N9
dffeas \rfile[27][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][21] .is_wysiwyg = "true";
defparam \rfile[27][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y28_N15
dffeas \rfile[31][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][21] .is_wysiwyg = "true";
defparam \rfile[31][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N31
dffeas \rfile[19][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][21] .is_wysiwyg = "true";
defparam \rfile[19][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N29
dffeas \rfile[23][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][21] .is_wysiwyg = "true";
defparam \rfile[23][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N30
cycloneive_lcell_comb \Mux42~7 (
// Equation(s):
// \Mux42~7_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[23][21]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[19][21]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[19][21]~q ),
	.datad(\rfile[23][21]~q ),
	.cin(gnd),
	.combout(\Mux42~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~7 .lut_mask = 16'hBA98;
defparam \Mux42~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N14
cycloneive_lcell_comb \Mux42~8 (
// Equation(s):
// \Mux42~8_combout  = (instruction_D[19] & ((\Mux42~7_combout  & ((\rfile[31][21]~q ))) # (!\Mux42~7_combout  & (\rfile[27][21]~q )))) # (!instruction_D[19] & (((\Mux42~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[27][21]~q ),
	.datac(\rfile[31][21]~q ),
	.datad(\Mux42~7_combout ),
	.cin(gnd),
	.combout(\Mux42~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~8 .lut_mask = 16'hF588;
defparam \Mux42~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y33_N13
dffeas \rfile[24][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][21] .is_wysiwyg = "true";
defparam \rfile[24][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y33_N7
dffeas \rfile[16][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][21] .is_wysiwyg = "true";
defparam \rfile[16][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N12
cycloneive_lcell_comb \Mux42~4 (
// Equation(s):
// \Mux42~4_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[24][21]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[16][21]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[24][21]~q ),
	.datad(\rfile[16][21]~q ),
	.cin(gnd),
	.combout(\Mux42~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~4 .lut_mask = 16'hB9A8;
defparam \Mux42~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N21
dffeas \rfile[28][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][21] .is_wysiwyg = "true";
defparam \rfile[28][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N20
cycloneive_lcell_comb \Mux42~5 (
// Equation(s):
// \Mux42~5_combout  = (\Mux42~4_combout  & (((\rfile[28][21]~q ) # (!instruction_D[18])))) # (!\Mux42~4_combout  & (\rfile[20][21]~q  & ((instruction_D[18]))))

	.dataa(\rfile[20][21]~q ),
	.datab(\Mux42~4_combout ),
	.datac(\rfile[28][21]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux42~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~5 .lut_mask = 16'hE2CC;
defparam \Mux42~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N3
dffeas \rfile[30][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][21] .is_wysiwyg = "true";
defparam \rfile[30][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y34_N17
dffeas \rfile[22][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][21] .is_wysiwyg = "true";
defparam \rfile[22][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N14
cycloneive_lcell_comb \rfile[26][21]~feeder (
// Equation(s):
// \rfile[26][21]~feeder_combout  = \wdat_WB[21]~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_21),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[26][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[26][21]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[26][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y36_N15
dffeas \rfile[26][21] (
	.clk(!CLK),
	.d(\rfile[26][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][21] .is_wysiwyg = "true";
defparam \rfile[26][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N12
cycloneive_lcell_comb \rfile[18][21]~feeder (
// Equation(s):
// \rfile[18][21]~feeder_combout  = \wdat_WB[21]~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_21),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[18][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[18][21]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[18][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N13
dffeas \rfile[18][21] (
	.clk(!CLK),
	.d(\rfile[18][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][21] .is_wysiwyg = "true";
defparam \rfile[18][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N0
cycloneive_lcell_comb \Mux42~2 (
// Equation(s):
// \Mux42~2_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[26][21]~q )) # (!instruction_D[19] & ((\rfile[18][21]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[26][21]~q ),
	.datad(\rfile[18][21]~q ),
	.cin(gnd),
	.combout(\Mux42~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~2 .lut_mask = 16'hD9C8;
defparam \Mux42~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N16
cycloneive_lcell_comb \Mux42~3 (
// Equation(s):
// \Mux42~3_combout  = (instruction_D[18] & ((\Mux42~2_combout  & (\rfile[30][21]~q )) # (!\Mux42~2_combout  & ((\rfile[22][21]~q ))))) # (!instruction_D[18] & (((\Mux42~2_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[30][21]~q ),
	.datac(\rfile[22][21]~q ),
	.datad(\Mux42~2_combout ),
	.cin(gnd),
	.combout(\Mux42~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~3 .lut_mask = 16'hDDA0;
defparam \Mux42~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N28
cycloneive_lcell_comb \Mux42~6 (
// Equation(s):
// \Mux42~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\Mux42~3_combout ))) # (!instruction_D[17] & (\Mux42~5_combout ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux42~5_combout ),
	.datad(\Mux42~3_combout ),
	.cin(gnd),
	.combout(\Mux42~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~6 .lut_mask = 16'hDC98;
defparam \Mux42~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N12
cycloneive_lcell_comb \rfile[14][21]~feeder (
// Equation(s):
// \rfile[14][21]~feeder_combout  = \wdat_WB[21]~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_21),
	.cin(gnd),
	.combout(\rfile[14][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][21]~feeder .lut_mask = 16'hFF00;
defparam \rfile[14][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N13
dffeas \rfile[14][21] (
	.clk(!CLK),
	.d(\rfile[14][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][21] .is_wysiwyg = "true";
defparam \rfile[14][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N31
dffeas \rfile[13][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][21] .is_wysiwyg = "true";
defparam \rfile[13][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N31
dffeas \rfile[12][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][21] .is_wysiwyg = "true";
defparam \rfile[12][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N30
cycloneive_lcell_comb \Mux42~17 (
// Equation(s):
// \Mux42~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][21]~q )))) # (!instruction_D[16] & (!instruction_D[17] & ((\rfile[12][21]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[13][21]~q ),
	.datad(\rfile[12][21]~q ),
	.cin(gnd),
	.combout(\Mux42~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~17 .lut_mask = 16'hB9A8;
defparam \Mux42~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N11
dffeas \rfile[15][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][21] .is_wysiwyg = "true";
defparam \rfile[15][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N12
cycloneive_lcell_comb \Mux42~18 (
// Equation(s):
// \Mux42~18_combout  = (instruction_D[17] & ((\Mux42~17_combout  & ((\rfile[15][21]~q ))) # (!\Mux42~17_combout  & (\rfile[14][21]~q )))) # (!instruction_D[17] & (((\Mux42~17_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[14][21]~q ),
	.datac(\Mux42~17_combout ),
	.datad(\rfile[15][21]~q ),
	.cin(gnd),
	.combout(\Mux42~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~18 .lut_mask = 16'hF858;
defparam \Mux42~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N16
cycloneive_lcell_comb \rfile[9][21]~feeder (
// Equation(s):
// \rfile[9][21]~feeder_combout  = \wdat_WB[21]~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_21),
	.cin(gnd),
	.combout(\rfile[9][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][21]~feeder .lut_mask = 16'hFF00;
defparam \rfile[9][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N17
dffeas \rfile[9][21] (
	.clk(!CLK),
	.d(\rfile[9][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][21] .is_wysiwyg = "true";
defparam \rfile[9][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N14
cycloneive_lcell_comb \rfile[11][21]~feeder (
// Equation(s):
// \rfile[11][21]~feeder_combout  = \wdat_WB[21]~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_21),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[11][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][21]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[11][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N15
dffeas \rfile[11][21] (
	.clk(!CLK),
	.d(\rfile[11][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][21] .is_wysiwyg = "true";
defparam \rfile[11][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N23
dffeas \rfile[8][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][21] .is_wysiwyg = "true";
defparam \rfile[8][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N1
dffeas \rfile[10][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][21] .is_wysiwyg = "true";
defparam \rfile[10][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N22
cycloneive_lcell_comb \Mux42~10 (
// Equation(s):
// \Mux42~10_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][21]~q ))) # (!instruction_D[17] & (\rfile[8][21]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[8][21]~q ),
	.datad(\rfile[10][21]~q ),
	.cin(gnd),
	.combout(\Mux42~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~10 .lut_mask = 16'hDC98;
defparam \Mux42~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N4
cycloneive_lcell_comb \Mux42~11 (
// Equation(s):
// \Mux42~11_combout  = (instruction_D[16] & ((\Mux42~10_combout  & ((\rfile[11][21]~q ))) # (!\Mux42~10_combout  & (\rfile[9][21]~q )))) # (!instruction_D[16] & (((\Mux42~10_combout ))))

	.dataa(\rfile[9][21]~q ),
	.datab(\rfile[11][21]~q ),
	.datac(instruction_D_16),
	.datad(\Mux42~10_combout ),
	.cin(gnd),
	.combout(\Mux42~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~11 .lut_mask = 16'hCFA0;
defparam \Mux42~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N27
dffeas \rfile[7][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][21] .is_wysiwyg = "true";
defparam \rfile[7][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N11
dffeas \rfile[6][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][21] .is_wysiwyg = "true";
defparam \rfile[6][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N29
dffeas \rfile[5][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][21] .is_wysiwyg = "true";
defparam \rfile[5][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N28
cycloneive_lcell_comb \Mux42~12 (
// Equation(s):
// \Mux42~12_combout  = (instruction_D[16] & (((\rfile[5][21]~q ) # (instruction_D[17])))) # (!instruction_D[16] & (\rfile[4][21]~q  & ((!instruction_D[17]))))

	.dataa(\rfile[4][21]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[5][21]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux42~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~12 .lut_mask = 16'hCCE2;
defparam \Mux42~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N10
cycloneive_lcell_comb \Mux42~13 (
// Equation(s):
// \Mux42~13_combout  = (instruction_D[17] & ((\Mux42~12_combout  & (\rfile[7][21]~q )) # (!\Mux42~12_combout  & ((\rfile[6][21]~q ))))) # (!instruction_D[17] & (((\Mux42~12_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[7][21]~q ),
	.datac(\rfile[6][21]~q ),
	.datad(\Mux42~12_combout ),
	.cin(gnd),
	.combout(\Mux42~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~13 .lut_mask = 16'hDDA0;
defparam \Mux42~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N11
dffeas \rfile[2][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][21] .is_wysiwyg = "true";
defparam \rfile[2][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N17
dffeas \rfile[3][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][21] .is_wysiwyg = "true";
defparam \rfile[3][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N11
dffeas \rfile[1][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][21] .is_wysiwyg = "true";
defparam \rfile[1][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N16
cycloneive_lcell_comb \Mux42~14 (
// Equation(s):
// \Mux42~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][21]~q )) # (!instruction_D[17] & ((\rfile[1][21]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[3][21]~q ),
	.datad(\rfile[1][21]~q ),
	.cin(gnd),
	.combout(\Mux42~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~14 .lut_mask = 16'hC480;
defparam \Mux42~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N28
cycloneive_lcell_comb \Mux42~15 (
// Equation(s):
// \Mux42~15_combout  = (\Mux42~14_combout ) # ((instruction_D[17] & (\rfile[2][21]~q  & !instruction_D[16])))

	.dataa(instruction_D_17),
	.datab(\rfile[2][21]~q ),
	.datac(instruction_D_16),
	.datad(\Mux42~14_combout ),
	.cin(gnd),
	.combout(\Mux42~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~15 .lut_mask = 16'hFF08;
defparam \Mux42~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N6
cycloneive_lcell_comb \Mux42~16 (
// Equation(s):
// \Mux42~16_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\Mux42~13_combout )))) # (!instruction_D[18] & (!instruction_D[19] & ((\Mux42~15_combout ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\Mux42~13_combout ),
	.datad(\Mux42~15_combout ),
	.cin(gnd),
	.combout(\Mux42~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~16 .lut_mask = 16'hB9A8;
defparam \Mux42~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N27
dffeas \rfile[29][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][20] .is_wysiwyg = "true";
defparam \rfile[29][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N9
dffeas \rfile[17][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][20] .is_wysiwyg = "true";
defparam \rfile[17][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N8
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[25][20]~q )) # (!instruction_D[19] & ((\rfile[17][20]~q )))))

	.dataa(\rfile[25][20]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[17][20]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hEE30;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N26
cycloneive_lcell_comb \rfile[21][20]~feeder (
// Equation(s):
// \rfile[21][20]~feeder_combout  = \wdat_WB[20]~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_20),
	.cin(gnd),
	.combout(\rfile[21][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][20]~feeder .lut_mask = 16'hFF00;
defparam \rfile[21][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N27
dffeas \rfile[21][20] (
	.clk(!CLK),
	.d(\rfile[21][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][20] .is_wysiwyg = "true";
defparam \rfile[21][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N4
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (instruction_D[18] & ((\Mux43~0_combout  & (\rfile[29][20]~q )) # (!\Mux43~0_combout  & ((\rfile[21][20]~q ))))) # (!instruction_D[18] & (((\Mux43~0_combout ))))

	.dataa(\rfile[29][20]~q ),
	.datab(instruction_D_18),
	.datac(\Mux43~0_combout ),
	.datad(\rfile[21][20]~q ),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hBCB0;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N19
dffeas \rfile[28][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][20] .is_wysiwyg = "true";
defparam \rfile[28][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y33_N26
cycloneive_lcell_comb \rfile[16][20]~feeder (
// Equation(s):
// \rfile[16][20]~feeder_combout  = \wdat_WB[20]~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_20),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[16][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[16][20]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[16][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y33_N27
dffeas \rfile[16][20] (
	.clk(!CLK),
	.d(\rfile[16][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][20] .is_wysiwyg = "true";
defparam \rfile[16][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y33_N0
cycloneive_lcell_comb \rfile[20][20]~feeder (
// Equation(s):
// \rfile[20][20]~feeder_combout  = \wdat_WB[20]~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_20),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[20][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[20][20]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[20][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y33_N1
dffeas \rfile[20][20] (
	.clk(!CLK),
	.d(\rfile[20][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][20] .is_wysiwyg = "true";
defparam \rfile[20][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y33_N24
cycloneive_lcell_comb \Mux43~4 (
// Equation(s):
// \Mux43~4_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[20][20]~q ))) # (!instruction_D[18] & (\rfile[16][20]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[16][20]~q ),
	.datad(\rfile[20][20]~q ),
	.cin(gnd),
	.combout(\Mux43~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~4 .lut_mask = 16'hDC98;
defparam \Mux43~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N18
cycloneive_lcell_comb \Mux43~5 (
// Equation(s):
// \Mux43~5_combout  = (instruction_D[19] & ((\Mux43~4_combout  & ((\rfile[28][20]~q ))) # (!\Mux43~4_combout  & (\rfile[24][20]~q )))) # (!instruction_D[19] & (((\Mux43~4_combout ))))

	.dataa(\rfile[24][20]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[28][20]~q ),
	.datad(\Mux43~4_combout ),
	.cin(gnd),
	.combout(\Mux43~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~5 .lut_mask = 16'hF388;
defparam \Mux43~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y34_N17
dffeas \rfile[30][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][20] .is_wysiwyg = "true";
defparam \rfile[30][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y34_N15
dffeas \rfile[26][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][20] .is_wysiwyg = "true";
defparam \rfile[26][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y35_N29
dffeas \rfile[18][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][20] .is_wysiwyg = "true";
defparam \rfile[18][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N28
cycloneive_lcell_comb \Mux43~2 (
// Equation(s):
// \Mux43~2_combout  = (instruction_D[18] & ((\rfile[22][20]~q ) # ((instruction_D[19])))) # (!instruction_D[18] & (((\rfile[18][20]~q  & !instruction_D[19]))))

	.dataa(\rfile[22][20]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[18][20]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux43~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~2 .lut_mask = 16'hCCB8;
defparam \Mux43~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N14
cycloneive_lcell_comb \Mux43~3 (
// Equation(s):
// \Mux43~3_combout  = (instruction_D[19] & ((\Mux43~2_combout  & (\rfile[30][20]~q )) # (!\Mux43~2_combout  & ((\rfile[26][20]~q ))))) # (!instruction_D[19] & (((\Mux43~2_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[30][20]~q ),
	.datac(\rfile[26][20]~q ),
	.datad(\Mux43~2_combout ),
	.cin(gnd),
	.combout(\Mux43~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~3 .lut_mask = 16'hDDA0;
defparam \Mux43~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N22
cycloneive_lcell_comb \Mux43~6 (
// Equation(s):
// \Mux43~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux43~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & (\Mux43~5_combout )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux43~5_combout ),
	.datad(\Mux43~3_combout ),
	.cin(gnd),
	.combout(\Mux43~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~6 .lut_mask = 16'hBA98;
defparam \Mux43~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y29_N21
dffeas \rfile[23][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][20] .is_wysiwyg = "true";
defparam \rfile[23][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N11
dffeas \rfile[19][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][20] .is_wysiwyg = "true";
defparam \rfile[19][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N29
dffeas \rfile[27][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][20] .is_wysiwyg = "true";
defparam \rfile[27][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N10
cycloneive_lcell_comb \Mux43~7 (
// Equation(s):
// \Mux43~7_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[27][20]~q )))) # (!instruction_D[19] & (!instruction_D[18] & (\rfile[19][20]~q )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[19][20]~q ),
	.datad(\rfile[27][20]~q ),
	.cin(gnd),
	.combout(\Mux43~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~7 .lut_mask = 16'hBA98;
defparam \Mux43~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N17
dffeas \rfile[31][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][20] .is_wysiwyg = "true";
defparam \rfile[31][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N16
cycloneive_lcell_comb \Mux43~8 (
// Equation(s):
// \Mux43~8_combout  = (\Mux43~7_combout  & (((\rfile[31][20]~q ) # (!instruction_D[18])))) # (!\Mux43~7_combout  & (\rfile[23][20]~q  & ((instruction_D[18]))))

	.dataa(\rfile[23][20]~q ),
	.datab(\Mux43~7_combout ),
	.datac(\rfile[31][20]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux43~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~8 .lut_mask = 16'hE2CC;
defparam \Mux43~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N1
dffeas \rfile[12][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][20] .is_wysiwyg = "true";
defparam \rfile[12][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N0
cycloneive_lcell_comb \rfile[13][20]~feeder (
// Equation(s):
// \rfile[13][20]~feeder_combout  = \wdat_WB[20]~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_20),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[13][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[13][20]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[13][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N1
dffeas \rfile[13][20] (
	.clk(!CLK),
	.d(\rfile[13][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][20] .is_wysiwyg = "true";
defparam \rfile[13][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N0
cycloneive_lcell_comb \Mux43~17 (
// Equation(s):
// \Mux43~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][20]~q ))) # (!instruction_D[16] & (\rfile[12][20]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][20]~q ),
	.datad(\rfile[13][20]~q ),
	.cin(gnd),
	.combout(\Mux43~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~17 .lut_mask = 16'hDC98;
defparam \Mux43~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N19
dffeas \rfile[14][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][20] .is_wysiwyg = "true";
defparam \rfile[14][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N9
dffeas \rfile[15][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][20] .is_wysiwyg = "true";
defparam \rfile[15][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N8
cycloneive_lcell_comb \Mux43~18 (
// Equation(s):
// \Mux43~18_combout  = (\Mux43~17_combout  & (((\rfile[15][20]~q ) # (!instruction_D[17])))) # (!\Mux43~17_combout  & (\rfile[14][20]~q  & ((instruction_D[17]))))

	.dataa(\Mux43~17_combout ),
	.datab(\rfile[14][20]~q ),
	.datac(\rfile[15][20]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux43~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~18 .lut_mask = 16'hE4AA;
defparam \Mux43~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N31
dffeas \rfile[2][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][20] .is_wysiwyg = "true";
defparam \rfile[2][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N1
dffeas \rfile[3][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][20] .is_wysiwyg = "true";
defparam \rfile[3][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N0
cycloneive_lcell_comb \Mux43~14 (
// Equation(s):
// \Mux43~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][20]~q ))) # (!instruction_D[17] & (\rfile[1][20]~q ))))

	.dataa(\rfile[1][20]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[3][20]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux43~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~14 .lut_mask = 16'hC088;
defparam \Mux43~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N30
cycloneive_lcell_comb \Mux43~15 (
// Equation(s):
// \Mux43~15_combout  = (\Mux43~14_combout ) # ((instruction_D[17] & (!instruction_D[16] & \rfile[2][20]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[2][20]~q ),
	.datad(\Mux43~14_combout ),
	.cin(gnd),
	.combout(\Mux43~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~15 .lut_mask = 16'hFF20;
defparam \Mux43~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N14
cycloneive_lcell_comb \rfile[9][20]~feeder (
// Equation(s):
// \rfile[9][20]~feeder_combout  = \wdat_WB[20]~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_20),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[9][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][20]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[9][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N15
dffeas \rfile[9][20] (
	.clk(!CLK),
	.d(\rfile[9][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][20] .is_wysiwyg = "true";
defparam \rfile[9][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N27
dffeas \rfile[8][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][20] .is_wysiwyg = "true";
defparam \rfile[8][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N17
dffeas \rfile[10][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][20] .is_wysiwyg = "true";
defparam \rfile[10][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N26
cycloneive_lcell_comb \Mux43~12 (
// Equation(s):
// \Mux43~12_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][20]~q )))) # (!instruction_D[17] & (!instruction_D[16] & (\rfile[8][20]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[8][20]~q ),
	.datad(\rfile[10][20]~q ),
	.cin(gnd),
	.combout(\Mux43~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~12 .lut_mask = 16'hBA98;
defparam \Mux43~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N20
cycloneive_lcell_comb \Mux43~13 (
// Equation(s):
// \Mux43~13_combout  = (instruction_D[16] & ((\Mux43~12_combout  & (\rfile[11][20]~q )) # (!\Mux43~12_combout  & ((\rfile[9][20]~q ))))) # (!instruction_D[16] & (((\Mux43~12_combout ))))

	.dataa(\rfile[11][20]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[9][20]~q ),
	.datad(\Mux43~12_combout ),
	.cin(gnd),
	.combout(\Mux43~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~13 .lut_mask = 16'hBBC0;
defparam \Mux43~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N24
cycloneive_lcell_comb \Mux43~16 (
// Equation(s):
// \Mux43~16_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\Mux43~13_combout )))) # (!instruction_D[19] & (!instruction_D[18] & (\Mux43~15_combout )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux43~15_combout ),
	.datad(\Mux43~13_combout ),
	.cin(gnd),
	.combout(\Mux43~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~16 .lut_mask = 16'hBA98;
defparam \Mux43~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y27_N7
dffeas \rfile[7][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][20] .is_wysiwyg = "true";
defparam \rfile[7][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N17
dffeas \rfile[4][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][20] .is_wysiwyg = "true";
defparam \rfile[4][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N11
dffeas \rfile[5][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][20] .is_wysiwyg = "true";
defparam \rfile[5][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N16
cycloneive_lcell_comb \Mux43~10 (
// Equation(s):
// \Mux43~10_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][20]~q ))) # (!instruction_D[16] & (\rfile[4][20]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][20]~q ),
	.datad(\rfile[5][20]~q ),
	.cin(gnd),
	.combout(\Mux43~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~10 .lut_mask = 16'hDC98;
defparam \Mux43~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N0
cycloneive_lcell_comb \rfile[6][20]~feeder (
// Equation(s):
// \rfile[6][20]~feeder_combout  = \wdat_WB[20]~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_20),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[6][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][20]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[6][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y27_N1
dffeas \rfile[6][20] (
	.clk(!CLK),
	.d(\rfile[6][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][20] .is_wysiwyg = "true";
defparam \rfile[6][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N16
cycloneive_lcell_comb \Mux43~11 (
// Equation(s):
// \Mux43~11_combout  = (instruction_D[17] & ((\Mux43~10_combout  & (\rfile[7][20]~q )) # (!\Mux43~10_combout  & ((\rfile[6][20]~q ))))) # (!instruction_D[17] & (((\Mux43~10_combout ))))

	.dataa(\rfile[7][20]~q ),
	.datab(instruction_D_17),
	.datac(\Mux43~10_combout ),
	.datad(\rfile[6][20]~q ),
	.cin(gnd),
	.combout(\Mux43~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~11 .lut_mask = 16'hBCB0;
defparam \Mux43~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N13
dffeas \rfile[29][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][19] .is_wysiwyg = "true";
defparam \rfile[29][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N11
dffeas \rfile[25][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][19] .is_wysiwyg = "true";
defparam \rfile[25][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N15
dffeas \rfile[21][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][19] .is_wysiwyg = "true";
defparam \rfile[21][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N23
dffeas \rfile[17][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][19] .is_wysiwyg = "true";
defparam \rfile[17][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N14
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[21][19]~q )) # (!instruction_D[18] & ((\rfile[17][19]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[21][19]~q ),
	.datad(\rfile[17][19]~q ),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hD9C8;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N10
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (instruction_D[19] & ((\Mux44~0_combout  & (\rfile[29][19]~q )) # (!\Mux44~0_combout  & ((\rfile[25][19]~q ))))) # (!instruction_D[19] & (((\Mux44~0_combout ))))

	.dataa(\rfile[29][19]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[25][19]~q ),
	.datad(\Mux44~0_combout ),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hBBC0;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y29_N19
dffeas \rfile[23][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][19] .is_wysiwyg = "true";
defparam \rfile[23][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N13
dffeas \rfile[19][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][19] .is_wysiwyg = "true";
defparam \rfile[19][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N18
cycloneive_lcell_comb \Mux44~7 (
// Equation(s):
// \Mux44~7_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[23][19]~q )) # (!instruction_D[18] & ((\rfile[19][19]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[23][19]~q ),
	.datad(\rfile[19][19]~q ),
	.cin(gnd),
	.combout(\Mux44~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~7 .lut_mask = 16'hD9C8;
defparam \Mux44~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N13
dffeas \rfile[31][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][19] .is_wysiwyg = "true";
defparam \rfile[31][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y29_N11
dffeas \rfile[27][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][19] .is_wysiwyg = "true";
defparam \rfile[27][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N12
cycloneive_lcell_comb \Mux44~8 (
// Equation(s):
// \Mux44~8_combout  = (instruction_D[19] & ((\Mux44~7_combout  & (\rfile[31][19]~q )) # (!\Mux44~7_combout  & ((\rfile[27][19]~q ))))) # (!instruction_D[19] & (\Mux44~7_combout ))

	.dataa(instruction_D_19),
	.datab(\Mux44~7_combout ),
	.datac(\rfile[31][19]~q ),
	.datad(\rfile[27][19]~q ),
	.cin(gnd),
	.combout(\Mux44~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~8 .lut_mask = 16'hE6C4;
defparam \Mux44~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N29
dffeas \rfile[20][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][19] .is_wysiwyg = "true";
defparam \rfile[20][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y33_N15
dffeas \rfile[28][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][19] .is_wysiwyg = "true";
defparam \rfile[28][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y33_N29
dffeas \rfile[16][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][19] .is_wysiwyg = "true";
defparam \rfile[16][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y33_N3
dffeas \rfile[24][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][19] .is_wysiwyg = "true";
defparam \rfile[24][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N28
cycloneive_lcell_comb \Mux44~4 (
// Equation(s):
// \Mux44~4_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[24][19]~q )))) # (!instruction_D[19] & (!instruction_D[18] & (\rfile[16][19]~q )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[16][19]~q ),
	.datad(\rfile[24][19]~q ),
	.cin(gnd),
	.combout(\Mux44~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~4 .lut_mask = 16'hBA98;
defparam \Mux44~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N14
cycloneive_lcell_comb \Mux44~5 (
// Equation(s):
// \Mux44~5_combout  = (instruction_D[18] & ((\Mux44~4_combout  & ((\rfile[28][19]~q ))) # (!\Mux44~4_combout  & (\rfile[20][19]~q )))) # (!instruction_D[18] & (((\Mux44~4_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[20][19]~q ),
	.datac(\rfile[28][19]~q ),
	.datad(\Mux44~4_combout ),
	.cin(gnd),
	.combout(\Mux44~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~5 .lut_mask = 16'hF588;
defparam \Mux44~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N15
dffeas \rfile[30][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][19] .is_wysiwyg = "true";
defparam \rfile[30][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y34_N25
dffeas \rfile[22][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][19] .is_wysiwyg = "true";
defparam \rfile[22][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y36_N23
dffeas \rfile[26][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][19] .is_wysiwyg = "true";
defparam \rfile[26][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N30
cycloneive_lcell_comb \rfile[18][19]~feeder (
// Equation(s):
// \rfile[18][19]~feeder_combout  = \wdat_WB[19]~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_19),
	.cin(gnd),
	.combout(\rfile[18][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[18][19]~feeder .lut_mask = 16'hFF00;
defparam \rfile[18][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N31
dffeas \rfile[18][19] (
	.clk(!CLK),
	.d(\rfile[18][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][19] .is_wysiwyg = "true";
defparam \rfile[18][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N22
cycloneive_lcell_comb \Mux44~2 (
// Equation(s):
// \Mux44~2_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[26][19]~q )) # (!instruction_D[19] & ((\rfile[18][19]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[26][19]~q ),
	.datad(\rfile[18][19]~q ),
	.cin(gnd),
	.combout(\Mux44~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~2 .lut_mask = 16'hD9C8;
defparam \Mux44~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N24
cycloneive_lcell_comb \Mux44~3 (
// Equation(s):
// \Mux44~3_combout  = (instruction_D[18] & ((\Mux44~2_combout  & (\rfile[30][19]~q )) # (!\Mux44~2_combout  & ((\rfile[22][19]~q ))))) # (!instruction_D[18] & (((\Mux44~2_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[30][19]~q ),
	.datac(\rfile[22][19]~q ),
	.datad(\Mux44~2_combout ),
	.cin(gnd),
	.combout(\Mux44~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~3 .lut_mask = 16'hDDA0;
defparam \Mux44~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N18
cycloneive_lcell_comb \Mux44~6 (
// Equation(s):
// \Mux44~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux44~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & (\Mux44~5_combout )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux44~5_combout ),
	.datad(\Mux44~3_combout ),
	.cin(gnd),
	.combout(\Mux44~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~6 .lut_mask = 16'hBA98;
defparam \Mux44~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y35_N7
dffeas \rfile[8][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][19] .is_wysiwyg = "true";
defparam \rfile[8][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N13
dffeas \rfile[10][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][19] .is_wysiwyg = "true";
defparam \rfile[10][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N6
cycloneive_lcell_comb \Mux44~10 (
// Equation(s):
// \Mux44~10_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][19]~q )))) # (!instruction_D[17] & (!instruction_D[16] & (\rfile[8][19]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[8][19]~q ),
	.datad(\rfile[10][19]~q ),
	.cin(gnd),
	.combout(\Mux44~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~10 .lut_mask = 16'hBA98;
defparam \Mux44~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N13
dffeas \rfile[11][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][19] .is_wysiwyg = "true";
defparam \rfile[11][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N19
dffeas \rfile[9][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][19] .is_wysiwyg = "true";
defparam \rfile[9][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N12
cycloneive_lcell_comb \Mux44~11 (
// Equation(s):
// \Mux44~11_combout  = (\Mux44~10_combout  & (((\rfile[11][19]~q )) # (!instruction_D[16]))) # (!\Mux44~10_combout  & (instruction_D[16] & ((\rfile[9][19]~q ))))

	.dataa(\Mux44~10_combout ),
	.datab(instruction_D_16),
	.datac(\rfile[11][19]~q ),
	.datad(\rfile[9][19]~q ),
	.cin(gnd),
	.combout(\Mux44~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~11 .lut_mask = 16'hE6A2;
defparam \Mux44~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N9
dffeas \rfile[6][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][19] .is_wysiwyg = "true";
defparam \rfile[6][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N3
dffeas \rfile[7][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][19] .is_wysiwyg = "true";
defparam \rfile[7][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N8
cycloneive_lcell_comb \Mux44~13 (
// Equation(s):
// \Mux44~13_combout  = (\Mux44~12_combout  & (((\rfile[7][19]~q )) # (!instruction_D[17]))) # (!\Mux44~12_combout  & (instruction_D[17] & (\rfile[6][19]~q )))

	.dataa(\Mux44~12_combout ),
	.datab(instruction_D_17),
	.datac(\rfile[6][19]~q ),
	.datad(\rfile[7][19]~q ),
	.cin(gnd),
	.combout(\Mux44~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~13 .lut_mask = 16'hEA62;
defparam \Mux44~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N7
dffeas \rfile[1][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][19] .is_wysiwyg = "true";
defparam \rfile[1][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N25
dffeas \rfile[3][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][19] .is_wysiwyg = "true";
defparam \rfile[3][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N6
cycloneive_lcell_comb \Mux44~14 (
// Equation(s):
// \Mux44~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][19]~q ))) # (!instruction_D[17] & (\rfile[1][19]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[1][19]~q ),
	.datad(\rfile[3][19]~q ),
	.cin(gnd),
	.combout(\Mux44~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~14 .lut_mask = 16'hC840;
defparam \Mux44~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N3
dffeas \rfile[2][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][19] .is_wysiwyg = "true";
defparam \rfile[2][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N0
cycloneive_lcell_comb \Mux44~15 (
// Equation(s):
// \Mux44~15_combout  = (\Mux44~14_combout ) # ((instruction_D[17] & (!instruction_D[16] & \rfile[2][19]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux44~14_combout ),
	.datad(\rfile[2][19]~q ),
	.cin(gnd),
	.combout(\Mux44~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~15 .lut_mask = 16'hF2F0;
defparam \Mux44~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N26
cycloneive_lcell_comb \Mux44~16 (
// Equation(s):
// \Mux44~16_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\Mux44~13_combout )) # (!instruction_D[18] & ((\Mux44~15_combout )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux44~13_combout ),
	.datad(\Mux44~15_combout ),
	.cin(gnd),
	.combout(\Mux44~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~16 .lut_mask = 16'hD9C8;
defparam \Mux44~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N16
cycloneive_lcell_comb \rfile[14][19]~feeder (
// Equation(s):
// \rfile[14][19]~feeder_combout  = \wdat_WB[19]~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_19),
	.cin(gnd),
	.combout(\rfile[14][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][19]~feeder .lut_mask = 16'hFF00;
defparam \rfile[14][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N17
dffeas \rfile[14][19] (
	.clk(!CLK),
	.d(\rfile[14][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][19] .is_wysiwyg = "true";
defparam \rfile[14][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N27
dffeas \rfile[15][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][19] .is_wysiwyg = "true";
defparam \rfile[15][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N25
dffeas \rfile[13][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][19] .is_wysiwyg = "true";
defparam \rfile[13][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N11
dffeas \rfile[12][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][19] .is_wysiwyg = "true";
defparam \rfile[12][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N24
cycloneive_lcell_comb \Mux44~17 (
// Equation(s):
// \Mux44~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[13][19]~q )) # (!instruction_D[16] & ((\rfile[12][19]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[13][19]~q ),
	.datad(\rfile[12][19]~q ),
	.cin(gnd),
	.combout(\Mux44~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~17 .lut_mask = 16'hD9C8;
defparam \Mux44~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N24
cycloneive_lcell_comb \Mux44~18 (
// Equation(s):
// \Mux44~18_combout  = (instruction_D[17] & ((\Mux44~17_combout  & ((\rfile[15][19]~q ))) # (!\Mux44~17_combout  & (\rfile[14][19]~q )))) # (!instruction_D[17] & (((\Mux44~17_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[14][19]~q ),
	.datac(\rfile[15][19]~q ),
	.datad(\Mux44~17_combout ),
	.cin(gnd),
	.combout(\Mux44~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~18 .lut_mask = 16'hF588;
defparam \Mux44~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N22
cycloneive_lcell_comb \rfile[21][18]~feeder (
// Equation(s):
// \rfile[21][18]~feeder_combout  = \wdat_WB[18]~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_18),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[21][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][18]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[21][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N23
dffeas \rfile[21][18] (
	.clk(!CLK),
	.d(\rfile[21][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][18] .is_wysiwyg = "true";
defparam \rfile[21][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N5
dffeas \rfile[29][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][18] .is_wysiwyg = "true";
defparam \rfile[29][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y30_N25
dffeas \rfile[17][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][18] .is_wysiwyg = "true";
defparam \rfile[17][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y30_N13
dffeas \rfile[25][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][18] .is_wysiwyg = "true";
defparam \rfile[25][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N24
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[25][18]~q ))) # (!instruction_D[19] & (\rfile[17][18]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[17][18]~q ),
	.datad(\rfile[25][18]~q ),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hDC98;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N4
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (instruction_D[18] & ((\Mux45~0_combout  & ((\rfile[29][18]~q ))) # (!\Mux45~0_combout  & (\rfile[21][18]~q )))) # (!instruction_D[18] & (((\Mux45~0_combout ))))

	.dataa(\rfile[21][18]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[29][18]~q ),
	.datad(\Mux45~0_combout ),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hF388;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N6
cycloneive_lcell_comb \rfile[23][18]~feeder (
// Equation(s):
// \rfile[23][18]~feeder_combout  = \wdat_WB[18]~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_18),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[23][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[23][18]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[23][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y31_N7
dffeas \rfile[23][18] (
	.clk(!CLK),
	.d(\rfile[23][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][18] .is_wysiwyg = "true";
defparam \rfile[23][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N1
dffeas \rfile[31][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][18] .is_wysiwyg = "true";
defparam \rfile[31][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y29_N31
dffeas \rfile[27][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][18] .is_wysiwyg = "true";
defparam \rfile[27][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N4
cycloneive_lcell_comb \rfile[19][18]~feeder (
// Equation(s):
// \rfile[19][18]~feeder_combout  = \wdat_WB[18]~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_18),
	.cin(gnd),
	.combout(\rfile[19][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[19][18]~feeder .lut_mask = 16'hFF00;
defparam \rfile[19][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y28_N5
dffeas \rfile[19][18] (
	.clk(!CLK),
	.d(\rfile[19][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][18] .is_wysiwyg = "true";
defparam \rfile[19][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N30
cycloneive_lcell_comb \Mux45~7 (
// Equation(s):
// \Mux45~7_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[27][18]~q )) # (!instruction_D[19] & ((\rfile[19][18]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[27][18]~q ),
	.datad(\rfile[19][18]~q ),
	.cin(gnd),
	.combout(\Mux45~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~7 .lut_mask = 16'hD9C8;
defparam \Mux45~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N0
cycloneive_lcell_comb \Mux45~8 (
// Equation(s):
// \Mux45~8_combout  = (instruction_D[18] & ((\Mux45~7_combout  & ((\rfile[31][18]~q ))) # (!\Mux45~7_combout  & (\rfile[23][18]~q )))) # (!instruction_D[18] & (((\Mux45~7_combout ))))

	.dataa(\rfile[23][18]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[31][18]~q ),
	.datad(\Mux45~7_combout ),
	.cin(gnd),
	.combout(\Mux45~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~8 .lut_mask = 16'hF388;
defparam \Mux45~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y34_N5
dffeas \rfile[30][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][18] .is_wysiwyg = "true";
defparam \rfile[30][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y34_N31
dffeas \rfile[26][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][18] .is_wysiwyg = "true";
defparam \rfile[26][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y35_N9
dffeas \rfile[18][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][18] .is_wysiwyg = "true";
defparam \rfile[18][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N10
cycloneive_lcell_comb \rfile[22][18]~feeder (
// Equation(s):
// \rfile[22][18]~feeder_combout  = \wdat_WB[18]~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_18),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[22][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[22][18]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[22][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y35_N11
dffeas \rfile[22][18] (
	.clk(!CLK),
	.d(\rfile[22][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][18] .is_wysiwyg = "true";
defparam \rfile[22][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N8
cycloneive_lcell_comb \Mux45~2 (
// Equation(s):
// \Mux45~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[22][18]~q ))) # (!instruction_D[18] & (\rfile[18][18]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][18]~q ),
	.datad(\rfile[22][18]~q ),
	.cin(gnd),
	.combout(\Mux45~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~2 .lut_mask = 16'hDC98;
defparam \Mux45~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N30
cycloneive_lcell_comb \Mux45~3 (
// Equation(s):
// \Mux45~3_combout  = (instruction_D[19] & ((\Mux45~2_combout  & (\rfile[30][18]~q )) # (!\Mux45~2_combout  & ((\rfile[26][18]~q ))))) # (!instruction_D[19] & (((\Mux45~2_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[30][18]~q ),
	.datac(\rfile[26][18]~q ),
	.datad(\Mux45~2_combout ),
	.cin(gnd),
	.combout(\Mux45~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~3 .lut_mask = 16'hDDA0;
defparam \Mux45~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N11
dffeas \rfile[28][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][18] .is_wysiwyg = "true";
defparam \rfile[28][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y33_N23
dffeas \rfile[24][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][18] .is_wysiwyg = "true";
defparam \rfile[24][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y33_N17
dffeas \rfile[16][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][18] .is_wysiwyg = "true";
defparam \rfile[16][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y33_N13
dffeas \rfile[20][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][18] .is_wysiwyg = "true";
defparam \rfile[20][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N16
cycloneive_lcell_comb \Mux45~4 (
// Equation(s):
// \Mux45~4_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[20][18]~q ))) # (!instruction_D[18] & (\rfile[16][18]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[16][18]~q ),
	.datad(\rfile[20][18]~q ),
	.cin(gnd),
	.combout(\Mux45~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~4 .lut_mask = 16'hDC98;
defparam \Mux45~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N22
cycloneive_lcell_comb \Mux45~5 (
// Equation(s):
// \Mux45~5_combout  = (instruction_D[19] & ((\Mux45~4_combout  & (\rfile[28][18]~q )) # (!\Mux45~4_combout  & ((\rfile[24][18]~q ))))) # (!instruction_D[19] & (((\Mux45~4_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[28][18]~q ),
	.datac(\rfile[24][18]~q ),
	.datad(\Mux45~4_combout ),
	.cin(gnd),
	.combout(\Mux45~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~5 .lut_mask = 16'hDDA0;
defparam \Mux45~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N16
cycloneive_lcell_comb \Mux45~6 (
// Equation(s):
// \Mux45~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\Mux45~3_combout )) # (!instruction_D[17] & ((\Mux45~5_combout )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux45~3_combout ),
	.datad(\Mux45~5_combout ),
	.cin(gnd),
	.combout(\Mux45~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~6 .lut_mask = 16'hD9C8;
defparam \Mux45~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N5
dffeas \rfile[4][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][18] .is_wysiwyg = "true";
defparam \rfile[4][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N6
cycloneive_lcell_comb \Mux45~10 (
// Equation(s):
// \Mux45~10_combout  = (instruction_D[16] & ((\rfile[5][18]~q ) # ((instruction_D[17])))) # (!instruction_D[16] & (((\rfile[4][18]~q  & !instruction_D[17]))))

	.dataa(\rfile[5][18]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[4][18]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux45~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~10 .lut_mask = 16'hCCB8;
defparam \Mux45~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N29
dffeas \rfile[7][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][18] .is_wysiwyg = "true";
defparam \rfile[7][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N30
cycloneive_lcell_comb \rfile[6][18]~feeder (
// Equation(s):
// \rfile[6][18]~feeder_combout  = \wdat_WB[18]~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_18),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[6][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][18]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[6][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N31
dffeas \rfile[6][18] (
	.clk(!CLK),
	.d(\rfile[6][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][18] .is_wysiwyg = "true";
defparam \rfile[6][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N28
cycloneive_lcell_comb \Mux45~11 (
// Equation(s):
// \Mux45~11_combout  = (\Mux45~10_combout  & (((\rfile[7][18]~q )) # (!instruction_D[17]))) # (!\Mux45~10_combout  & (instruction_D[17] & ((\rfile[6][18]~q ))))

	.dataa(\Mux45~10_combout ),
	.datab(instruction_D_17),
	.datac(\rfile[7][18]~q ),
	.datad(\rfile[6][18]~q ),
	.cin(gnd),
	.combout(\Mux45~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~11 .lut_mask = 16'hE6A2;
defparam \Mux45~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N5
dffeas \rfile[15][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][18] .is_wysiwyg = "true";
defparam \rfile[15][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N11
dffeas \rfile[14][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][18] .is_wysiwyg = "true";
defparam \rfile[14][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N1
dffeas \rfile[13][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][18] .is_wysiwyg = "true";
defparam \rfile[13][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N7
dffeas \rfile[12][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][18] .is_wysiwyg = "true";
defparam \rfile[12][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N0
cycloneive_lcell_comb \Mux45~17 (
// Equation(s):
// \Mux45~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[13][18]~q )) # (!instruction_D[16] & ((\rfile[12][18]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[13][18]~q ),
	.datad(\rfile[12][18]~q ),
	.cin(gnd),
	.combout(\Mux45~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~17 .lut_mask = 16'hD9C8;
defparam \Mux45~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N10
cycloneive_lcell_comb \Mux45~18 (
// Equation(s):
// \Mux45~18_combout  = (instruction_D[17] & ((\Mux45~17_combout  & (\rfile[15][18]~q )) # (!\Mux45~17_combout  & ((\rfile[14][18]~q ))))) # (!instruction_D[17] & (((\Mux45~17_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[15][18]~q ),
	.datac(\rfile[14][18]~q ),
	.datad(\Mux45~17_combout ),
	.cin(gnd),
	.combout(\Mux45~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~18 .lut_mask = 16'hDDA0;
defparam \Mux45~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N9
dffeas \rfile[2][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][18] .is_wysiwyg = "true";
defparam \rfile[2][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y31_N15
dffeas \rfile[1][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][18] .is_wysiwyg = "true";
defparam \rfile[1][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N0
cycloneive_lcell_comb \rfile[3][18]~feeder (
// Equation(s):
// \rfile[3][18]~feeder_combout  = \wdat_WB[18]~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_18),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[3][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[3][18]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[3][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N1
dffeas \rfile[3][18] (
	.clk(!CLK),
	.d(\rfile[3][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][18] .is_wysiwyg = "true";
defparam \rfile[3][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N12
cycloneive_lcell_comb \Mux45~14 (
// Equation(s):
// \Mux45~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][18]~q ))) # (!instruction_D[17] & (\rfile[1][18]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[1][18]~q ),
	.datad(\rfile[3][18]~q ),
	.cin(gnd),
	.combout(\Mux45~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~14 .lut_mask = 16'hA820;
defparam \Mux45~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N8
cycloneive_lcell_comb \Mux45~15 (
// Equation(s):
// \Mux45~15_combout  = (\Mux45~14_combout ) # ((!instruction_D[16] & (instruction_D[17] & \rfile[2][18]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[2][18]~q ),
	.datad(\Mux45~14_combout ),
	.cin(gnd),
	.combout(\Mux45~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~15 .lut_mask = 16'hFF40;
defparam \Mux45~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N16
cycloneive_lcell_comb \rfile[11][18]~feeder (
// Equation(s):
// \rfile[11][18]~feeder_combout  = \wdat_WB[18]~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_18),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[11][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][18]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[11][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N17
dffeas \rfile[11][18] (
	.clk(!CLK),
	.d(\rfile[11][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][18] .is_wysiwyg = "true";
defparam \rfile[11][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N15
dffeas \rfile[9][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][18] .is_wysiwyg = "true";
defparam \rfile[9][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N5
dffeas \rfile[8][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][18] .is_wysiwyg = "true";
defparam \rfile[8][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N6
cycloneive_lcell_comb \rfile[10][18]~feeder (
// Equation(s):
// \rfile[10][18]~feeder_combout  = \wdat_WB[18]~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_18),
	.cin(gnd),
	.combout(\rfile[10][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[10][18]~feeder .lut_mask = 16'hFF00;
defparam \rfile[10][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N7
dffeas \rfile[10][18] (
	.clk(!CLK),
	.d(\rfile[10][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][18] .is_wysiwyg = "true";
defparam \rfile[10][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N4
cycloneive_lcell_comb \Mux45~12 (
// Equation(s):
// \Mux45~12_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][18]~q ))) # (!instruction_D[17] & (\rfile[8][18]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[8][18]~q ),
	.datad(\rfile[10][18]~q ),
	.cin(gnd),
	.combout(\Mux45~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~12 .lut_mask = 16'hDC98;
defparam \Mux45~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N14
cycloneive_lcell_comb \Mux45~13 (
// Equation(s):
// \Mux45~13_combout  = (instruction_D[16] & ((\Mux45~12_combout  & (\rfile[11][18]~q )) # (!\Mux45~12_combout  & ((\rfile[9][18]~q ))))) # (!instruction_D[16] & (((\Mux45~12_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][18]~q ),
	.datac(\rfile[9][18]~q ),
	.datad(\Mux45~12_combout ),
	.cin(gnd),
	.combout(\Mux45~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~13 .lut_mask = 16'hDDA0;
defparam \Mux45~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N2
cycloneive_lcell_comb \Mux45~16 (
// Equation(s):
// \Mux45~16_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\Mux45~13_combout )))) # (!instruction_D[19] & (!instruction_D[18] & (\Mux45~15_combout )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux45~15_combout ),
	.datad(\Mux45~13_combout ),
	.cin(gnd),
	.combout(\Mux45~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~16 .lut_mask = 16'hBA98;
defparam \Mux45~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N15
dffeas \rfile[28][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][17] .is_wysiwyg = "true";
defparam \rfile[28][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y33_N15
dffeas \rfile[24][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][17] .is_wysiwyg = "true";
defparam \rfile[24][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y33_N1
dffeas \rfile[16][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][17] .is_wysiwyg = "true";
defparam \rfile[16][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N14
cycloneive_lcell_comb \Mux46~4 (
// Equation(s):
// \Mux46~4_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[24][17]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[16][17]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[24][17]~q ),
	.datad(\rfile[16][17]~q ),
	.cin(gnd),
	.combout(\Mux46~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~4 .lut_mask = 16'hB9A8;
defparam \Mux46~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N8
cycloneive_lcell_comb \Mux46~5 (
// Equation(s):
// \Mux46~5_combout  = (instruction_D[18] & ((\Mux46~4_combout  & ((\rfile[28][17]~q ))) # (!\Mux46~4_combout  & (\rfile[20][17]~q )))) # (!instruction_D[18] & (((\Mux46~4_combout ))))

	.dataa(\rfile[20][17]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[28][17]~q ),
	.datad(\Mux46~4_combout ),
	.cin(gnd),
	.combout(\Mux46~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~5 .lut_mask = 16'hF388;
defparam \Mux46~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y35_N17
dffeas \rfile[30][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][17] .is_wysiwyg = "true";
defparam \rfile[30][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N15
dffeas \rfile[18][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][17] .is_wysiwyg = "true";
defparam \rfile[18][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N29
dffeas \rfile[26][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][17] .is_wysiwyg = "true";
defparam \rfile[26][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N28
cycloneive_lcell_comb \Mux46~2 (
// Equation(s):
// \Mux46~2_combout  = (instruction_D[19] & (((\rfile[26][17]~q ) # (instruction_D[18])))) # (!instruction_D[19] & (\rfile[18][17]~q  & ((!instruction_D[18]))))

	.dataa(instruction_D_19),
	.datab(\rfile[18][17]~q ),
	.datac(\rfile[26][17]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~2 .lut_mask = 16'hAAE4;
defparam \Mux46~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N16
cycloneive_lcell_comb \Mux46~3 (
// Equation(s):
// \Mux46~3_combout  = (instruction_D[18] & ((\Mux46~2_combout  & ((\rfile[30][17]~q ))) # (!\Mux46~2_combout  & (\rfile[22][17]~q )))) # (!instruction_D[18] & (((\Mux46~2_combout ))))

	.dataa(\rfile[22][17]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[30][17]~q ),
	.datad(\Mux46~2_combout ),
	.cin(gnd),
	.combout(\Mux46~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~3 .lut_mask = 16'hF388;
defparam \Mux46~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N2
cycloneive_lcell_comb \Mux46~6 (
// Equation(s):
// \Mux46~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux46~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & (\Mux46~5_combout )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux46~5_combout ),
	.datad(\Mux46~3_combout ),
	.cin(gnd),
	.combout(\Mux46~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~6 .lut_mask = 16'hBA98;
defparam \Mux46~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y28_N0
cycloneive_lcell_comb \rfile[27][17]~feeder (
// Equation(s):
// \rfile[27][17]~feeder_combout  = \wdat_WB[17]~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_17),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[27][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[27][17]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[27][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y28_N1
dffeas \rfile[27][17] (
	.clk(!CLK),
	.d(\rfile[27][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][17] .is_wysiwyg = "true";
defparam \rfile[27][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y28_N17
dffeas \rfile[31][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][17] .is_wysiwyg = "true";
defparam \rfile[31][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N15
dffeas \rfile[23][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][17] .is_wysiwyg = "true";
defparam \rfile[23][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N30
cycloneive_lcell_comb \rfile[19][17]~feeder (
// Equation(s):
// \rfile[19][17]~feeder_combout  = \wdat_WB[17]~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_17),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[19][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[19][17]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[19][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y28_N31
dffeas \rfile[19][17] (
	.clk(!CLK),
	.d(\rfile[19][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][17] .is_wysiwyg = "true";
defparam \rfile[19][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N14
cycloneive_lcell_comb \Mux46~7 (
// Equation(s):
// \Mux46~7_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[23][17]~q )) # (!instruction_D[18] & ((\rfile[19][17]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[23][17]~q ),
	.datad(\rfile[19][17]~q ),
	.cin(gnd),
	.combout(\Mux46~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~7 .lut_mask = 16'hD9C8;
defparam \Mux46~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N16
cycloneive_lcell_comb \Mux46~8 (
// Equation(s):
// \Mux46~8_combout  = (instruction_D[19] & ((\Mux46~7_combout  & ((\rfile[31][17]~q ))) # (!\Mux46~7_combout  & (\rfile[27][17]~q )))) # (!instruction_D[19] & (((\Mux46~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[27][17]~q ),
	.datac(\rfile[31][17]~q ),
	.datad(\Mux46~7_combout ),
	.cin(gnd),
	.combout(\Mux46~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~8 .lut_mask = 16'hF588;
defparam \Mux46~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N25
dffeas \rfile[29][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][17] .is_wysiwyg = "true";
defparam \rfile[29][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N31
dffeas \rfile[25][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][17] .is_wysiwyg = "true";
defparam \rfile[25][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y30_N23
dffeas \rfile[17][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][17] .is_wysiwyg = "true";
defparam \rfile[17][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N0
cycloneive_lcell_comb \rfile[21][17]~feeder (
// Equation(s):
// \rfile[21][17]~feeder_combout  = \wdat_WB[17]~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_17),
	.cin(gnd),
	.combout(\rfile[21][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][17]~feeder .lut_mask = 16'hFF00;
defparam \rfile[21][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y28_N1
dffeas \rfile[21][17] (
	.clk(!CLK),
	.d(\rfile[21][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][17] .is_wysiwyg = "true";
defparam \rfile[21][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N22
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[21][17]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[17][17]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[17][17]~q ),
	.datad(\rfile[21][17]~q ),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hBA98;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N30
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (instruction_D[19] & ((\Mux46~0_combout  & (\rfile[29][17]~q )) # (!\Mux46~0_combout  & ((\rfile[25][17]~q ))))) # (!instruction_D[19] & (((\Mux46~0_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[29][17]~q ),
	.datac(\rfile[25][17]~q ),
	.datad(\Mux46~0_combout ),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hDDA0;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N8
cycloneive_lcell_comb \rfile[6][17]~feeder (
// Equation(s):
// \rfile[6][17]~feeder_combout  = \wdat_WB[17]~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_17),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[6][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][17]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[6][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N9
dffeas \rfile[6][17] (
	.clk(!CLK),
	.d(\rfile[6][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][17] .is_wysiwyg = "true";
defparam \rfile[6][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N29
dffeas \rfile[7][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][17] .is_wysiwyg = "true";
defparam \rfile[7][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N5
dffeas \rfile[5][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][17] .is_wysiwyg = "true";
defparam \rfile[5][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N23
dffeas \rfile[4][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][17] .is_wysiwyg = "true";
defparam \rfile[4][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N22
cycloneive_lcell_comb \Mux46~12 (
// Equation(s):
// \Mux46~12_combout  = (instruction_D[16] & ((\rfile[5][17]~q ) # ((instruction_D[17])))) # (!instruction_D[16] & (((\rfile[4][17]~q  & !instruction_D[17]))))

	.dataa(instruction_D_16),
	.datab(\rfile[5][17]~q ),
	.datac(\rfile[4][17]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux46~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~12 .lut_mask = 16'hAAD8;
defparam \Mux46~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N10
cycloneive_lcell_comb \Mux46~13 (
// Equation(s):
// \Mux46~13_combout  = (instruction_D[17] & ((\Mux46~12_combout  & ((\rfile[7][17]~q ))) # (!\Mux46~12_combout  & (\rfile[6][17]~q )))) # (!instruction_D[17] & (((\Mux46~12_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[6][17]~q ),
	.datac(\rfile[7][17]~q ),
	.datad(\Mux46~12_combout ),
	.cin(gnd),
	.combout(\Mux46~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~13 .lut_mask = 16'hF588;
defparam \Mux46~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N31
dffeas \rfile[3][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][17] .is_wysiwyg = "true";
defparam \rfile[3][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y31_N29
dffeas \rfile[1][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][17] .is_wysiwyg = "true";
defparam \rfile[1][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N30
cycloneive_lcell_comb \Mux46~14 (
// Equation(s):
// \Mux46~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][17]~q )) # (!instruction_D[17] & ((\rfile[1][17]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[3][17]~q ),
	.datad(\rfile[1][17]~q ),
	.cin(gnd),
	.combout(\Mux46~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~14 .lut_mask = 16'hA280;
defparam \Mux46~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N0
cycloneive_lcell_comb \rfile[2][17]~feeder (
// Equation(s):
// \rfile[2][17]~feeder_combout  = \wdat_WB[17]~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_17),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[2][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][17]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[2][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N1
dffeas \rfile[2][17] (
	.clk(!CLK),
	.d(\rfile[2][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][17] .is_wysiwyg = "true";
defparam \rfile[2][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N22
cycloneive_lcell_comb \Mux46~15 (
// Equation(s):
// \Mux46~15_combout  = (\Mux46~14_combout ) # ((!instruction_D[16] & (instruction_D[17] & \rfile[2][17]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux46~14_combout ),
	.datad(\rfile[2][17]~q ),
	.cin(gnd),
	.combout(\Mux46~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~15 .lut_mask = 16'hF4F0;
defparam \Mux46~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N4
cycloneive_lcell_comb \Mux46~16 (
// Equation(s):
// \Mux46~16_combout  = (instruction_D[18] & ((\Mux46~13_combout ) # ((instruction_D[19])))) # (!instruction_D[18] & (((\Mux46~15_combout  & !instruction_D[19]))))

	.dataa(\Mux46~13_combout ),
	.datab(instruction_D_18),
	.datac(\Mux46~15_combout ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux46~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~16 .lut_mask = 16'hCCB8;
defparam \Mux46~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N1
dffeas \rfile[9][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][17] .is_wysiwyg = "true";
defparam \rfile[9][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N31
dffeas \rfile[11][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][17] .is_wysiwyg = "true";
defparam \rfile[11][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N21
dffeas \rfile[10][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][17] .is_wysiwyg = "true";
defparam \rfile[10][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N3
dffeas \rfile[8][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][17] .is_wysiwyg = "true";
defparam \rfile[8][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N20
cycloneive_lcell_comb \Mux46~10 (
// Equation(s):
// \Mux46~10_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][17]~q )))) # (!instruction_D[17] & (!instruction_D[16] & ((\rfile[8][17]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[10][17]~q ),
	.datad(\rfile[8][17]~q ),
	.cin(gnd),
	.combout(\Mux46~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~10 .lut_mask = 16'hB9A8;
defparam \Mux46~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N30
cycloneive_lcell_comb \Mux46~11 (
// Equation(s):
// \Mux46~11_combout  = (instruction_D[16] & ((\Mux46~10_combout  & ((\rfile[11][17]~q ))) # (!\Mux46~10_combout  & (\rfile[9][17]~q )))) # (!instruction_D[16] & (((\Mux46~10_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[9][17]~q ),
	.datac(\rfile[11][17]~q ),
	.datad(\Mux46~10_combout ),
	.cin(gnd),
	.combout(\Mux46~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~11 .lut_mask = 16'hF588;
defparam \Mux46~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N29
dffeas \rfile[15][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][17] .is_wysiwyg = "true";
defparam \rfile[15][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N27
dffeas \rfile[14][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][17] .is_wysiwyg = "true";
defparam \rfile[14][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N31
dffeas \rfile[12][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][17] .is_wysiwyg = "true";
defparam \rfile[12][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N26
cycloneive_lcell_comb \rfile[13][17]~feeder (
// Equation(s):
// \rfile[13][17]~feeder_combout  = \wdat_WB[17]~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_17),
	.cin(gnd),
	.combout(\rfile[13][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[13][17]~feeder .lut_mask = 16'hFF00;
defparam \rfile[13][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N27
dffeas \rfile[13][17] (
	.clk(!CLK),
	.d(\rfile[13][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][17] .is_wysiwyg = "true";
defparam \rfile[13][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N30
cycloneive_lcell_comb \Mux46~17 (
// Equation(s):
// \Mux46~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][17]~q ))) # (!instruction_D[16] & (\rfile[12][17]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][17]~q ),
	.datad(\rfile[13][17]~q ),
	.cin(gnd),
	.combout(\Mux46~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~17 .lut_mask = 16'hDC98;
defparam \Mux46~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N26
cycloneive_lcell_comb \Mux46~18 (
// Equation(s):
// \Mux46~18_combout  = (instruction_D[17] & ((\Mux46~17_combout  & (\rfile[15][17]~q )) # (!\Mux46~17_combout  & ((\rfile[14][17]~q ))))) # (!instruction_D[17] & (((\Mux46~17_combout ))))

	.dataa(\rfile[15][17]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[14][17]~q ),
	.datad(\Mux46~17_combout ),
	.cin(gnd),
	.combout(\Mux46~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~18 .lut_mask = 16'hBBC0;
defparam \Mux46~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y29_N27
dffeas \rfile[19][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][16] .is_wysiwyg = "true";
defparam \rfile[19][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N13
dffeas \rfile[27][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][16] .is_wysiwyg = "true";
defparam \rfile[27][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N26
cycloneive_lcell_comb \Mux47~7 (
// Equation(s):
// \Mux47~7_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[27][16]~q )))) # (!instruction_D[19] & (!instruction_D[18] & (\rfile[19][16]~q )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[19][16]~q ),
	.datad(\rfile[27][16]~q ),
	.cin(gnd),
	.combout(\Mux47~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~7 .lut_mask = 16'hBA98;
defparam \Mux47~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y29_N9
dffeas \rfile[23][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][16] .is_wysiwyg = "true";
defparam \rfile[23][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y29_N7
dffeas \rfile[31][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][16] .is_wysiwyg = "true";
defparam \rfile[31][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N8
cycloneive_lcell_comb \Mux47~8 (
// Equation(s):
// \Mux47~8_combout  = (\Mux47~7_combout  & (((\rfile[31][16]~q )) # (!instruction_D[18]))) # (!\Mux47~7_combout  & (instruction_D[18] & (\rfile[23][16]~q )))

	.dataa(\Mux47~7_combout ),
	.datab(instruction_D_18),
	.datac(\rfile[23][16]~q ),
	.datad(\rfile[31][16]~q ),
	.cin(gnd),
	.combout(\Mux47~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~8 .lut_mask = 16'hEA62;
defparam \Mux47~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y30_N5
dffeas \rfile[28][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][16] .is_wysiwyg = "true";
defparam \rfile[28][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N8
cycloneive_lcell_comb \rfile[20][16]~feeder (
// Equation(s):
// \rfile[20][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_16),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[20][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[20][16]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[20][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y30_N9
dffeas \rfile[20][16] (
	.clk(!CLK),
	.d(\rfile[20][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][16] .is_wysiwyg = "true";
defparam \rfile[20][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N18
cycloneive_lcell_comb \rfile[16][16]~feeder (
// Equation(s):
// \rfile[16][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_16),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[16][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[16][16]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[16][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y30_N19
dffeas \rfile[16][16] (
	.clk(!CLK),
	.d(\rfile[16][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][16] .is_wysiwyg = "true";
defparam \rfile[16][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N16
cycloneive_lcell_comb \Mux47~4 (
// Equation(s):
// \Mux47~4_combout  = (instruction_D[18] & ((\rfile[20][16]~q ) # ((instruction_D[19])))) # (!instruction_D[18] & (((!instruction_D[19] & \rfile[16][16]~q ))))

	.dataa(instruction_D_18),
	.datab(\rfile[20][16]~q ),
	.datac(instruction_D_19),
	.datad(\rfile[16][16]~q ),
	.cin(gnd),
	.combout(\Mux47~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~4 .lut_mask = 16'hADA8;
defparam \Mux47~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N4
cycloneive_lcell_comb \Mux47~5 (
// Equation(s):
// \Mux47~5_combout  = (instruction_D[19] & ((\Mux47~4_combout  & ((\rfile[28][16]~q ))) # (!\Mux47~4_combout  & (\rfile[24][16]~q )))) # (!instruction_D[19] & (((\Mux47~4_combout ))))

	.dataa(\rfile[24][16]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[28][16]~q ),
	.datad(\Mux47~4_combout ),
	.cin(gnd),
	.combout(\Mux47~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~5 .lut_mask = 16'hF388;
defparam \Mux47~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y35_N13
dffeas \rfile[30][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][16] .is_wysiwyg = "true";
defparam \rfile[30][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N5
dffeas \rfile[26][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][16] .is_wysiwyg = "true";
defparam \rfile[26][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N4
cycloneive_lcell_comb \Mux47~3 (
// Equation(s):
// \Mux47~3_combout  = (\Mux47~2_combout  & ((\rfile[30][16]~q ) # ((!instruction_D[19])))) # (!\Mux47~2_combout  & (((\rfile[26][16]~q  & instruction_D[19]))))

	.dataa(\Mux47~2_combout ),
	.datab(\rfile[30][16]~q ),
	.datac(\rfile[26][16]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux47~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~3 .lut_mask = 16'hD8AA;
defparam \Mux47~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N8
cycloneive_lcell_comb \Mux47~6 (
// Equation(s):
// \Mux47~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\Mux47~3_combout ))) # (!instruction_D[17] & (\Mux47~5_combout ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux47~5_combout ),
	.datad(\Mux47~3_combout ),
	.cin(gnd),
	.combout(\Mux47~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~6 .lut_mask = 16'hDC98;
defparam \Mux47~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N15
dffeas \rfile[29][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][16] .is_wysiwyg = "true";
defparam \rfile[29][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N12
cycloneive_lcell_comb \rfile[21][16]~feeder (
// Equation(s):
// \rfile[21][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_16),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[21][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][16]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[21][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N13
dffeas \rfile[21][16] (
	.clk(!CLK),
	.d(\rfile[21][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][16] .is_wysiwyg = "true";
defparam \rfile[21][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y30_N29
dffeas \rfile[17][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][16] .is_wysiwyg = "true";
defparam \rfile[17][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y30_N19
dffeas \rfile[25][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][16] .is_wysiwyg = "true";
defparam \rfile[25][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N28
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[25][16]~q ))) # (!instruction_D[19] & (\rfile[17][16]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[17][16]~q ),
	.datad(\rfile[25][16]~q ),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hDC98;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N2
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (instruction_D[18] & ((\Mux47~0_combout  & (\rfile[29][16]~q )) # (!\Mux47~0_combout  & ((\rfile[21][16]~q ))))) # (!instruction_D[18] & (((\Mux47~0_combout ))))

	.dataa(\rfile[29][16]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[21][16]~q ),
	.datad(\Mux47~0_combout ),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hBBC0;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N8
cycloneive_lcell_comb \rfile[9][16]~feeder (
// Equation(s):
// \rfile[9][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_16),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[9][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][16]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[9][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N9
dffeas \rfile[9][16] (
	.clk(!CLK),
	.d(\rfile[9][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][16] .is_wysiwyg = "true";
defparam \rfile[9][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y29_N17
dffeas \rfile[11][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][16] .is_wysiwyg = "true";
defparam \rfile[11][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N1
dffeas \rfile[10][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][16] .is_wysiwyg = "true";
defparam \rfile[10][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N0
cycloneive_lcell_comb \Mux47~12 (
// Equation(s):
// \Mux47~12_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][16]~q ))) # (!instruction_D[17] & (\rfile[8][16]~q ))))

	.dataa(\rfile[8][16]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[10][16]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux47~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~12 .lut_mask = 16'hFC22;
defparam \Mux47~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N18
cycloneive_lcell_comb \Mux47~13 (
// Equation(s):
// \Mux47~13_combout  = (instruction_D[16] & ((\Mux47~12_combout  & ((\rfile[11][16]~q ))) # (!\Mux47~12_combout  & (\rfile[9][16]~q )))) # (!instruction_D[16] & (((\Mux47~12_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[9][16]~q ),
	.datac(\rfile[11][16]~q ),
	.datad(\Mux47~12_combout ),
	.cin(gnd),
	.combout(\Mux47~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~13 .lut_mask = 16'hF588;
defparam \Mux47~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N31
dffeas \rfile[1][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][16] .is_wysiwyg = "true";
defparam \rfile[1][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N17
dffeas \rfile[3][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][16] .is_wysiwyg = "true";
defparam \rfile[3][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N30
cycloneive_lcell_comb \Mux47~14 (
// Equation(s):
// \Mux47~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][16]~q ))) # (!instruction_D[17] & (\rfile[1][16]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[1][16]~q ),
	.datad(\rfile[3][16]~q ),
	.cin(gnd),
	.combout(\Mux47~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~14 .lut_mask = 16'hC840;
defparam \Mux47~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N26
cycloneive_lcell_comb \rfile[2][16]~feeder (
// Equation(s):
// \rfile[2][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_16),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[2][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][16]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[2][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y29_N27
dffeas \rfile[2][16] (
	.clk(!CLK),
	.d(\rfile[2][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][16] .is_wysiwyg = "true";
defparam \rfile[2][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N20
cycloneive_lcell_comb \Mux47~15 (
// Equation(s):
// \Mux47~15_combout  = (\Mux47~14_combout ) # ((instruction_D[17] & (\rfile[2][16]~q  & !instruction_D[16])))

	.dataa(instruction_D_17),
	.datab(\Mux47~14_combout ),
	.datac(\rfile[2][16]~q ),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux47~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~15 .lut_mask = 16'hCCEC;
defparam \Mux47~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N22
cycloneive_lcell_comb \Mux47~16 (
// Equation(s):
// \Mux47~16_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\Mux47~13_combout )))) # (!instruction_D[19] & (!instruction_D[18] & ((\Mux47~15_combout ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux47~13_combout ),
	.datad(\Mux47~15_combout ),
	.cin(gnd),
	.combout(\Mux47~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~16 .lut_mask = 16'hB9A8;
defparam \Mux47~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N30
cycloneive_lcell_comb \rfile[6][16]~feeder (
// Equation(s):
// \rfile[6][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_16),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[6][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][16]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[6][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y27_N31
dffeas \rfile[6][16] (
	.clk(!CLK),
	.d(\rfile[6][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][16] .is_wysiwyg = "true";
defparam \rfile[6][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N21
dffeas \rfile[7][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][16] .is_wysiwyg = "true";
defparam \rfile[7][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N1
dffeas \rfile[5][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][16] .is_wysiwyg = "true";
defparam \rfile[5][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N0
cycloneive_lcell_comb \Mux47~10 (
// Equation(s):
// \Mux47~10_combout  = (instruction_D[16] & (((\rfile[5][16]~q ) # (instruction_D[17])))) # (!instruction_D[16] & (\rfile[4][16]~q  & ((!instruction_D[17]))))

	.dataa(\rfile[4][16]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[5][16]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux47~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~10 .lut_mask = 16'hCCE2;
defparam \Mux47~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N20
cycloneive_lcell_comb \Mux47~11 (
// Equation(s):
// \Mux47~11_combout  = (instruction_D[17] & ((\Mux47~10_combout  & ((\rfile[7][16]~q ))) # (!\Mux47~10_combout  & (\rfile[6][16]~q )))) # (!instruction_D[17] & (((\Mux47~10_combout ))))

	.dataa(\rfile[6][16]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[7][16]~q ),
	.datad(\Mux47~10_combout ),
	.cin(gnd),
	.combout(\Mux47~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~11 .lut_mask = 16'hF388;
defparam \Mux47~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N22
cycloneive_lcell_comb \rfile[14][16]~feeder (
// Equation(s):
// \rfile[14][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_16),
	.cin(gnd),
	.combout(\rfile[14][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][16]~feeder .lut_mask = 16'hFF00;
defparam \rfile[14][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N23
dffeas \rfile[14][16] (
	.clk(!CLK),
	.d(\rfile[14][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][16] .is_wysiwyg = "true";
defparam \rfile[14][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N0
cycloneive_lcell_comb \rfile[15][16]~feeder (
// Equation(s):
// \rfile[15][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_16),
	.cin(gnd),
	.combout(\rfile[15][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][16]~feeder .lut_mask = 16'hFF00;
defparam \rfile[15][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N1
dffeas \rfile[15][16] (
	.clk(!CLK),
	.d(\rfile[15][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][16] .is_wysiwyg = "true";
defparam \rfile[15][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N9
dffeas \rfile[12][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][16] .is_wysiwyg = "true";
defparam \rfile[12][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N24
cycloneive_lcell_comb \rfile[13][16]~feeder (
// Equation(s):
// \rfile[13][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_16),
	.cin(gnd),
	.combout(\rfile[13][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[13][16]~feeder .lut_mask = 16'hFF00;
defparam \rfile[13][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N25
dffeas \rfile[13][16] (
	.clk(!CLK),
	.d(\rfile[13][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][16] .is_wysiwyg = "true";
defparam \rfile[13][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N8
cycloneive_lcell_comb \Mux47~17 (
// Equation(s):
// \Mux47~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][16]~q ))) # (!instruction_D[16] & (\rfile[12][16]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][16]~q ),
	.datad(\rfile[13][16]~q ),
	.cin(gnd),
	.combout(\Mux47~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~17 .lut_mask = 16'hDC98;
defparam \Mux47~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N14
cycloneive_lcell_comb \Mux47~18 (
// Equation(s):
// \Mux47~18_combout  = (instruction_D[17] & ((\Mux47~17_combout  & ((\rfile[15][16]~q ))) # (!\Mux47~17_combout  & (\rfile[14][16]~q )))) # (!instruction_D[17] & (((\Mux47~17_combout ))))

	.dataa(\rfile[14][16]~q ),
	.datab(\rfile[15][16]~q ),
	.datac(instruction_D_17),
	.datad(\Mux47~17_combout ),
	.cin(gnd),
	.combout(\Mux47~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~18 .lut_mask = 16'hCFA0;
defparam \Mux47~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N29
dffeas \rfile[21][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][15] .is_wysiwyg = "true";
defparam \rfile[21][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N18
cycloneive_lcell_comb \rfile[17][15]~feeder (
// Equation(s):
// \rfile[17][15]~feeder_combout  = \wdat_WB[15]~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_15),
	.cin(gnd),
	.combout(\rfile[17][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[17][15]~feeder .lut_mask = 16'hFF00;
defparam \rfile[17][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N19
dffeas \rfile[17][15] (
	.clk(!CLK),
	.d(\rfile[17][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][15] .is_wysiwyg = "true";
defparam \rfile[17][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N26
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (instruction_D[18] & ((\rfile[21][15]~q ) # ((instruction_D[19])))) # (!instruction_D[18] & (((!instruction_D[19] & \rfile[17][15]~q ))))

	.dataa(instruction_D_18),
	.datab(\rfile[21][15]~q ),
	.datac(instruction_D_19),
	.datad(\rfile[17][15]~q ),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hADA8;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N5
dffeas \rfile[25][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][15] .is_wysiwyg = "true";
defparam \rfile[25][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N11
dffeas \rfile[29][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][15] .is_wysiwyg = "true";
defparam \rfile[29][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N4
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (\Mux48~0_combout  & (((\rfile[29][15]~q )) # (!instruction_D[19]))) # (!\Mux48~0_combout  & (instruction_D[19] & (\rfile[25][15]~q )))

	.dataa(\Mux48~0_combout ),
	.datab(instruction_D_19),
	.datac(\rfile[25][15]~q ),
	.datad(\rfile[29][15]~q ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'hEA62;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y29_N17
dffeas \rfile[27][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][15] .is_wysiwyg = "true";
defparam \rfile[27][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N3
dffeas \rfile[31][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][15] .is_wysiwyg = "true";
defparam \rfile[31][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N13
dffeas \rfile[23][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][15] .is_wysiwyg = "true";
defparam \rfile[23][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N3
dffeas \rfile[19][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][15] .is_wysiwyg = "true";
defparam \rfile[19][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N12
cycloneive_lcell_comb \Mux48~7 (
// Equation(s):
// \Mux48~7_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[23][15]~q )) # (!instruction_D[18] & ((\rfile[19][15]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[23][15]~q ),
	.datad(\rfile[19][15]~q ),
	.cin(gnd),
	.combout(\Mux48~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~7 .lut_mask = 16'hD9C8;
defparam \Mux48~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N2
cycloneive_lcell_comb \Mux48~8 (
// Equation(s):
// \Mux48~8_combout  = (instruction_D[19] & ((\Mux48~7_combout  & ((\rfile[31][15]~q ))) # (!\Mux48~7_combout  & (\rfile[27][15]~q )))) # (!instruction_D[19] & (((\Mux48~7_combout ))))

	.dataa(\rfile[27][15]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[31][15]~q ),
	.datad(\Mux48~7_combout ),
	.cin(gnd),
	.combout(\Mux48~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~8 .lut_mask = 16'hF388;
defparam \Mux48~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N24
cycloneive_lcell_comb \rfile[30][15]~feeder (
// Equation(s):
// \rfile[30][15]~feeder_combout  = \wdat_WB[15]~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_15),
	.cin(gnd),
	.combout(\rfile[30][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[30][15]~feeder .lut_mask = 16'hFF00;
defparam \rfile[30][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N25
dffeas \rfile[30][15] (
	.clk(!CLK),
	.d(\rfile[30][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][15] .is_wysiwyg = "true";
defparam \rfile[30][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y30_N1
dffeas \rfile[22][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][15] .is_wysiwyg = "true";
defparam \rfile[22][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N7
dffeas \rfile[18][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][15] .is_wysiwyg = "true";
defparam \rfile[18][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N21
dffeas \rfile[26][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][15] .is_wysiwyg = "true";
defparam \rfile[26][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N6
cycloneive_lcell_comb \Mux48~2 (
// Equation(s):
// \Mux48~2_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[26][15]~q ))) # (!instruction_D[19] & (\rfile[18][15]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[18][15]~q ),
	.datad(\rfile[26][15]~q ),
	.cin(gnd),
	.combout(\Mux48~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~2 .lut_mask = 16'hDC98;
defparam \Mux48~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N10
cycloneive_lcell_comb \Mux48~3 (
// Equation(s):
// \Mux48~3_combout  = (instruction_D[18] & ((\Mux48~2_combout  & (\rfile[30][15]~q )) # (!\Mux48~2_combout  & ((\rfile[22][15]~q ))))) # (!instruction_D[18] & (((\Mux48~2_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[30][15]~q ),
	.datac(\rfile[22][15]~q ),
	.datad(\Mux48~2_combout ),
	.cin(gnd),
	.combout(\Mux48~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~3 .lut_mask = 16'hDDA0;
defparam \Mux48~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y32_N27
dffeas \rfile[20][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][15] .is_wysiwyg = "true";
defparam \rfile[20][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y33_N21
dffeas \rfile[16][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][15] .is_wysiwyg = "true";
defparam \rfile[16][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N20
cycloneive_lcell_comb \Mux48~4 (
// Equation(s):
// \Mux48~4_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[24][15]~q )) # (!instruction_D[19] & ((\rfile[16][15]~q )))))

	.dataa(\rfile[24][15]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[16][15]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux48~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~4 .lut_mask = 16'hEE30;
defparam \Mux48~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N26
cycloneive_lcell_comb \Mux48~5 (
// Equation(s):
// \Mux48~5_combout  = (instruction_D[18] & ((\Mux48~4_combout  & (\rfile[28][15]~q )) # (!\Mux48~4_combout  & ((\rfile[20][15]~q ))))) # (!instruction_D[18] & (((\Mux48~4_combout ))))

	.dataa(\rfile[28][15]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[20][15]~q ),
	.datad(\Mux48~4_combout ),
	.cin(gnd),
	.combout(\Mux48~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~5 .lut_mask = 16'hBBC0;
defparam \Mux48~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N24
cycloneive_lcell_comb \Mux48~6 (
// Equation(s):
// \Mux48~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux48~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & ((\Mux48~5_combout ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux48~3_combout ),
	.datad(\Mux48~5_combout ),
	.cin(gnd),
	.combout(\Mux48~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~6 .lut_mask = 16'hB9A8;
defparam \Mux48~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N24
cycloneive_lcell_comb \rfile[14][15]~feeder (
// Equation(s):
// \rfile[14][15]~feeder_combout  = \wdat_WB[15]~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_15),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[14][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][15]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[14][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N25
dffeas \rfile[14][15] (
	.clk(!CLK),
	.d(\rfile[14][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][15] .is_wysiwyg = "true";
defparam \rfile[14][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N30
cycloneive_lcell_comb \rfile[15][15]~feeder (
// Equation(s):
// \rfile[15][15]~feeder_combout  = \wdat_WB[15]~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_15),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[15][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][15]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[15][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N31
dffeas \rfile[15][15] (
	.clk(!CLK),
	.d(\rfile[15][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][15] .is_wysiwyg = "true";
defparam \rfile[15][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N15
dffeas \rfile[12][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][15] .is_wysiwyg = "true";
defparam \rfile[12][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N9
dffeas \rfile[13][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][15] .is_wysiwyg = "true";
defparam \rfile[13][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N8
cycloneive_lcell_comb \Mux48~17 (
// Equation(s):
// \Mux48~17_combout  = (instruction_D[17] & (((instruction_D[16])))) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][15]~q ))) # (!instruction_D[16] & (\rfile[12][15]~q ))))

	.dataa(instruction_D_17),
	.datab(\rfile[12][15]~q ),
	.datac(\rfile[13][15]~q ),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux48~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~17 .lut_mask = 16'hFA44;
defparam \Mux48~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N14
cycloneive_lcell_comb \Mux48~18 (
// Equation(s):
// \Mux48~18_combout  = (instruction_D[17] & ((\Mux48~17_combout  & ((\rfile[15][15]~q ))) # (!\Mux48~17_combout  & (\rfile[14][15]~q )))) # (!instruction_D[17] & (((\Mux48~17_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[14][15]~q ),
	.datac(\rfile[15][15]~q ),
	.datad(\Mux48~17_combout ),
	.cin(gnd),
	.combout(\Mux48~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~18 .lut_mask = 16'hF588;
defparam \Mux48~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N27
dffeas \rfile[9][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][15] .is_wysiwyg = "true";
defparam \rfile[9][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y29_N9
dffeas \rfile[11][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][15] .is_wysiwyg = "true";
defparam \rfile[11][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N9
dffeas \rfile[10][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][15] .is_wysiwyg = "true";
defparam \rfile[10][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N31
dffeas \rfile[8][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][15] .is_wysiwyg = "true";
defparam \rfile[8][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N30
cycloneive_lcell_comb \Mux48~10 (
// Equation(s):
// \Mux48~10_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & (\rfile[10][15]~q )) # (!instruction_D[17] & ((\rfile[8][15]~q )))))

	.dataa(instruction_D_16),
	.datab(\rfile[10][15]~q ),
	.datac(\rfile[8][15]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux48~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~10 .lut_mask = 16'hEE50;
defparam \Mux48~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N22
cycloneive_lcell_comb \Mux48~11 (
// Equation(s):
// \Mux48~11_combout  = (\Mux48~10_combout  & (((\rfile[11][15]~q ) # (!instruction_D[16])))) # (!\Mux48~10_combout  & (\rfile[9][15]~q  & ((instruction_D[16]))))

	.dataa(\rfile[9][15]~q ),
	.datab(\rfile[11][15]~q ),
	.datac(\Mux48~10_combout ),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux48~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~11 .lut_mask = 16'hCAF0;
defparam \Mux48~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N0
cycloneive_lcell_comb \rfile[2][15]~feeder (
// Equation(s):
// \rfile[2][15]~feeder_combout  = \wdat_WB[15]~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_15),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[2][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][15]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[2][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y29_N1
dffeas \rfile[2][15] (
	.clk(!CLK),
	.d(\rfile[2][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][15] .is_wysiwyg = "true";
defparam \rfile[2][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N7
dffeas \rfile[3][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][15] .is_wysiwyg = "true";
defparam \rfile[3][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N25
dffeas \rfile[1][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][15] .is_wysiwyg = "true";
defparam \rfile[1][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N6
cycloneive_lcell_comb \Mux48~14 (
// Equation(s):
// \Mux48~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][15]~q )) # (!instruction_D[17] & ((\rfile[1][15]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[3][15]~q ),
	.datad(\rfile[1][15]~q ),
	.cin(gnd),
	.combout(\Mux48~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~14 .lut_mask = 16'hC480;
defparam \Mux48~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N6
cycloneive_lcell_comb \Mux48~15 (
// Equation(s):
// \Mux48~15_combout  = (\Mux48~14_combout ) # ((instruction_D[17] & (\rfile[2][15]~q  & !instruction_D[16])))

	.dataa(instruction_D_17),
	.datab(\rfile[2][15]~q ),
	.datac(\Mux48~14_combout ),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux48~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~15 .lut_mask = 16'hF0F8;
defparam \Mux48~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y27_N25
dffeas \rfile[7][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][15] .is_wysiwyg = "true";
defparam \rfile[7][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N27
dffeas \rfile[6][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][15] .is_wysiwyg = "true";
defparam \rfile[6][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N24
cycloneive_lcell_comb \rfile[5][15]~feeder (
// Equation(s):
// \rfile[5][15]~feeder_combout  = \wdat_WB[15]~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_15),
	.cin(gnd),
	.combout(\rfile[5][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[5][15]~feeder .lut_mask = 16'hFF00;
defparam \rfile[5][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N25
dffeas \rfile[5][15] (
	.clk(!CLK),
	.d(\rfile[5][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][15] .is_wysiwyg = "true";
defparam \rfile[5][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N20
cycloneive_lcell_comb \rfile[4][15]~feeder (
// Equation(s):
// \rfile[4][15]~feeder_combout  = \wdat_WB[15]~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_15),
	.cin(gnd),
	.combout(\rfile[4][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[4][15]~feeder .lut_mask = 16'hFF00;
defparam \rfile[4][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N21
dffeas \rfile[4][15] (
	.clk(!CLK),
	.d(\rfile[4][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][15] .is_wysiwyg = "true";
defparam \rfile[4][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N18
cycloneive_lcell_comb \Mux48~12 (
// Equation(s):
// \Mux48~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[5][15]~q )) # (!instruction_D[16] & ((\rfile[4][15]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[5][15]~q ),
	.datad(\rfile[4][15]~q ),
	.cin(gnd),
	.combout(\Mux48~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~12 .lut_mask = 16'hD9C8;
defparam \Mux48~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N26
cycloneive_lcell_comb \Mux48~13 (
// Equation(s):
// \Mux48~13_combout  = (instruction_D[17] & ((\Mux48~12_combout  & (\rfile[7][15]~q )) # (!\Mux48~12_combout  & ((\rfile[6][15]~q ))))) # (!instruction_D[17] & (((\Mux48~12_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[7][15]~q ),
	.datac(\rfile[6][15]~q ),
	.datad(\Mux48~12_combout ),
	.cin(gnd),
	.combout(\Mux48~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~13 .lut_mask = 16'hDDA0;
defparam \Mux48~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N20
cycloneive_lcell_comb \Mux48~16 (
// Equation(s):
// \Mux48~16_combout  = (instruction_D[19] & (((instruction_D[18])))) # (!instruction_D[19] & ((instruction_D[18] & ((\Mux48~13_combout ))) # (!instruction_D[18] & (\Mux48~15_combout ))))

	.dataa(\Mux48~15_combout ),
	.datab(instruction_D_19),
	.datac(instruction_D_18),
	.datad(\Mux48~13_combout ),
	.cin(gnd),
	.combout(\Mux48~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~16 .lut_mask = 16'hF2C2;
defparam \Mux48~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y29_N27
dffeas \rfile[31][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][14] .is_wysiwyg = "true";
defparam \rfile[31][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y29_N17
dffeas \rfile[23][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][14] .is_wysiwyg = "true";
defparam \rfile[23][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N15
dffeas \rfile[27][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][14] .is_wysiwyg = "true";
defparam \rfile[27][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N1
dffeas \rfile[19][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][14] .is_wysiwyg = "true";
defparam \rfile[19][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N0
cycloneive_lcell_comb \Mux49~7 (
// Equation(s):
// \Mux49~7_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[27][14]~q )) # (!instruction_D[19] & ((\rfile[19][14]~q )))))

	.dataa(instruction_D_18),
	.datab(\rfile[27][14]~q ),
	.datac(\rfile[19][14]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux49~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~7 .lut_mask = 16'hEE50;
defparam \Mux49~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N16
cycloneive_lcell_comb \Mux49~8 (
// Equation(s):
// \Mux49~8_combout  = (instruction_D[18] & ((\Mux49~7_combout  & (\rfile[31][14]~q )) # (!\Mux49~7_combout  & ((\rfile[23][14]~q ))))) # (!instruction_D[18] & (((\Mux49~7_combout ))))

	.dataa(\rfile[31][14]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[23][14]~q ),
	.datad(\Mux49~7_combout ),
	.cin(gnd),
	.combout(\Mux49~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~8 .lut_mask = 16'hBBC0;
defparam \Mux49~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y35_N9
dffeas \rfile[30][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][14] .is_wysiwyg = "true";
defparam \rfile[30][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N13
dffeas \rfile[26][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][14] .is_wysiwyg = "true";
defparam \rfile[26][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N3
dffeas \rfile[18][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][14] .is_wysiwyg = "true";
defparam \rfile[18][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y35_N19
dffeas \rfile[22][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][14] .is_wysiwyg = "true";
defparam \rfile[22][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N2
cycloneive_lcell_comb \Mux49~2 (
// Equation(s):
// \Mux49~2_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[22][14]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[18][14]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[18][14]~q ),
	.datad(\rfile[22][14]~q ),
	.cin(gnd),
	.combout(\Mux49~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~2 .lut_mask = 16'hBA98;
defparam \Mux49~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N12
cycloneive_lcell_comb \Mux49~3 (
// Equation(s):
// \Mux49~3_combout  = (instruction_D[19] & ((\Mux49~2_combout  & (\rfile[30][14]~q )) # (!\Mux49~2_combout  & ((\rfile[26][14]~q ))))) # (!instruction_D[19] & (((\Mux49~2_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[30][14]~q ),
	.datac(\rfile[26][14]~q ),
	.datad(\Mux49~2_combout ),
	.cin(gnd),
	.combout(\Mux49~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~3 .lut_mask = 16'hDDA0;
defparam \Mux49~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y30_N29
dffeas \rfile[28][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][14] .is_wysiwyg = "true";
defparam \rfile[28][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y32_N21
dffeas \rfile[20][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][14] .is_wysiwyg = "true";
defparam \rfile[20][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y32_N31
dffeas \rfile[16][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][14] .is_wysiwyg = "true";
defparam \rfile[16][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N30
cycloneive_lcell_comb \Mux49~4 (
// Equation(s):
// \Mux49~4_combout  = (instruction_D[19] & (((instruction_D[18])))) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[20][14]~q )) # (!instruction_D[18] & ((\rfile[16][14]~q )))))

	.dataa(instruction_D_19),
	.datab(\rfile[20][14]~q ),
	.datac(\rfile[16][14]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux49~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~4 .lut_mask = 16'hEE50;
defparam \Mux49~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N28
cycloneive_lcell_comb \Mux49~5 (
// Equation(s):
// \Mux49~5_combout  = (instruction_D[19] & ((\Mux49~4_combout  & ((\rfile[28][14]~q ))) # (!\Mux49~4_combout  & (\rfile[24][14]~q )))) # (!instruction_D[19] & (((\Mux49~4_combout ))))

	.dataa(\rfile[24][14]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[28][14]~q ),
	.datad(\Mux49~4_combout ),
	.cin(gnd),
	.combout(\Mux49~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~5 .lut_mask = 16'hF388;
defparam \Mux49~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N0
cycloneive_lcell_comb \Mux49~6 (
// Equation(s):
// \Mux49~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux49~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & ((\Mux49~5_combout ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux49~3_combout ),
	.datad(\Mux49~5_combout ),
	.cin(gnd),
	.combout(\Mux49~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~6 .lut_mask = 16'hB9A8;
defparam \Mux49~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N0
cycloneive_lcell_comb \rfile[21][14]~feeder (
// Equation(s):
// \rfile[21][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_14),
	.cin(gnd),
	.combout(\rfile[21][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][14]~feeder .lut_mask = 16'hFF00;
defparam \rfile[21][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N1
dffeas \rfile[21][14] (
	.clk(!CLK),
	.d(\rfile[21][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][14] .is_wysiwyg = "true";
defparam \rfile[21][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N18
cycloneive_lcell_comb \rfile[29][14]~feeder (
// Equation(s):
// \rfile[29][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_14),
	.cin(gnd),
	.combout(\rfile[29][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[29][14]~feeder .lut_mask = 16'hFF00;
defparam \rfile[29][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N19
dffeas \rfile[29][14] (
	.clk(!CLK),
	.d(\rfile[29][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][14] .is_wysiwyg = "true";
defparam \rfile[29][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y30_N21
dffeas \rfile[17][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][14] .is_wysiwyg = "true";
defparam \rfile[17][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N2
cycloneive_lcell_comb \rfile[25][14]~feeder (
// Equation(s):
// \rfile[25][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_14),
	.cin(gnd),
	.combout(\rfile[25][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[25][14]~feeder .lut_mask = 16'hFF00;
defparam \rfile[25][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N3
dffeas \rfile[25][14] (
	.clk(!CLK),
	.d(\rfile[25][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][14] .is_wysiwyg = "true";
defparam \rfile[25][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N20
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[25][14]~q ))) # (!instruction_D[19] & (\rfile[17][14]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[17][14]~q ),
	.datad(\rfile[25][14]~q ),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'hDC98;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N28
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (instruction_D[18] & ((\Mux49~0_combout  & ((\rfile[29][14]~q ))) # (!\Mux49~0_combout  & (\rfile[21][14]~q )))) # (!instruction_D[18] & (((\Mux49~0_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[21][14]~q ),
	.datac(\rfile[29][14]~q ),
	.datad(\Mux49~0_combout ),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hF588;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N16
cycloneive_lcell_comb \rfile[14][14]~feeder (
// Equation(s):
// \rfile[14][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_14),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[14][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][14]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[14][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N17
dffeas \rfile[14][14] (
	.clk(!CLK),
	.d(\rfile[14][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][14] .is_wysiwyg = "true";
defparam \rfile[14][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N10
cycloneive_lcell_comb \rfile[15][14]~feeder (
// Equation(s):
// \rfile[15][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_14),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[15][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][14]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[15][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N11
dffeas \rfile[15][14] (
	.clk(!CLK),
	.d(\rfile[15][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][14] .is_wysiwyg = "true";
defparam \rfile[15][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N19
dffeas \rfile[12][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][14] .is_wysiwyg = "true";
defparam \rfile[12][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N16
cycloneive_lcell_comb \rfile[13][14]~feeder (
// Equation(s):
// \rfile[13][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_14),
	.cin(gnd),
	.combout(\rfile[13][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[13][14]~feeder .lut_mask = 16'hFF00;
defparam \rfile[13][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N17
dffeas \rfile[13][14] (
	.clk(!CLK),
	.d(\rfile[13][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][14] .is_wysiwyg = "true";
defparam \rfile[13][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N18
cycloneive_lcell_comb \Mux49~17 (
// Equation(s):
// \Mux49~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][14]~q ))) # (!instruction_D[16] & (\rfile[12][14]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][14]~q ),
	.datad(\rfile[13][14]~q ),
	.cin(gnd),
	.combout(\Mux49~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~17 .lut_mask = 16'hDC98;
defparam \Mux49~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N6
cycloneive_lcell_comb \Mux49~18 (
// Equation(s):
// \Mux49~18_combout  = (instruction_D[17] & ((\Mux49~17_combout  & ((\rfile[15][14]~q ))) # (!\Mux49~17_combout  & (\rfile[14][14]~q )))) # (!instruction_D[17] & (((\Mux49~17_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[14][14]~q ),
	.datac(\rfile[15][14]~q ),
	.datad(\Mux49~17_combout ),
	.cin(gnd),
	.combout(\Mux49~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~18 .lut_mask = 16'hF588;
defparam \Mux49~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N2
cycloneive_lcell_comb \rfile[2][14]~feeder (
// Equation(s):
// \rfile[2][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_14),
	.cin(gnd),
	.combout(\rfile[2][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][14]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N3
dffeas \rfile[2][14] (
	.clk(!CLK),
	.d(\rfile[2][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][14] .is_wysiwyg = "true";
defparam \rfile[2][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y30_N29
dffeas \rfile[1][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][14] .is_wysiwyg = "true";
defparam \rfile[1][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y30_N3
dffeas \rfile[3][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][14] .is_wysiwyg = "true";
defparam \rfile[3][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N28
cycloneive_lcell_comb \Mux49~14 (
// Equation(s):
// \Mux49~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][14]~q ))) # (!instruction_D[17] & (\rfile[1][14]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[1][14]~q ),
	.datad(\rfile[3][14]~q ),
	.cin(gnd),
	.combout(\Mux49~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~14 .lut_mask = 16'hC840;
defparam \Mux49~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N14
cycloneive_lcell_comb \Mux49~15 (
// Equation(s):
// \Mux49~15_combout  = (\Mux49~14_combout ) # ((instruction_D[17] & (!instruction_D[16] & \rfile[2][14]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[2][14]~q ),
	.datad(\Mux49~14_combout ),
	.cin(gnd),
	.combout(\Mux49~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~15 .lut_mask = 16'hFF20;
defparam \Mux49~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N14
cycloneive_lcell_comb \rfile[11][14]~feeder (
// Equation(s):
// \rfile[11][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_14),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[11][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][14]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[11][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N15
dffeas \rfile[11][14] (
	.clk(!CLK),
	.d(\rfile[11][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][14] .is_wysiwyg = "true";
defparam \rfile[11][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N17
dffeas \rfile[9][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][14] .is_wysiwyg = "true";
defparam \rfile[9][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N17
dffeas \rfile[10][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][14] .is_wysiwyg = "true";
defparam \rfile[10][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N11
dffeas \rfile[8][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][14] .is_wysiwyg = "true";
defparam \rfile[8][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N16
cycloneive_lcell_comb \Mux49~12 (
// Equation(s):
// \Mux49~12_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\rfile[10][14]~q )) # (!instruction_D[17] & ((\rfile[8][14]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[10][14]~q ),
	.datad(\rfile[8][14]~q ),
	.cin(gnd),
	.combout(\Mux49~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~12 .lut_mask = 16'hD9C8;
defparam \Mux49~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N16
cycloneive_lcell_comb \Mux49~13 (
// Equation(s):
// \Mux49~13_combout  = (instruction_D[16] & ((\Mux49~12_combout  & (\rfile[11][14]~q )) # (!\Mux49~12_combout  & ((\rfile[9][14]~q ))))) # (!instruction_D[16] & (((\Mux49~12_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][14]~q ),
	.datac(\rfile[9][14]~q ),
	.datad(\Mux49~12_combout ),
	.cin(gnd),
	.combout(\Mux49~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~13 .lut_mask = 16'hDDA0;
defparam \Mux49~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N8
cycloneive_lcell_comb \Mux49~16 (
// Equation(s):
// \Mux49~16_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\Mux49~13_combout )))) # (!instruction_D[19] & (!instruction_D[18] & (\Mux49~15_combout )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux49~15_combout ),
	.datad(\Mux49~13_combout ),
	.cin(gnd),
	.combout(\Mux49~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~16 .lut_mask = 16'hBA98;
defparam \Mux49~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N22
cycloneive_lcell_comb \rfile[7][14]~feeder (
// Equation(s):
// \rfile[7][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_14),
	.cin(gnd),
	.combout(\rfile[7][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[7][14]~feeder .lut_mask = 16'hFF00;
defparam \rfile[7][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N23
dffeas \rfile[7][14] (
	.clk(!CLK),
	.d(\rfile[7][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][14] .is_wysiwyg = "true";
defparam \rfile[7][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N24
cycloneive_lcell_comb \rfile[6][14]~feeder (
// Equation(s):
// \rfile[6][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_14),
	.cin(gnd),
	.combout(\rfile[6][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][14]~feeder .lut_mask = 16'hFF00;
defparam \rfile[6][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N25
dffeas \rfile[6][14] (
	.clk(!CLK),
	.d(\rfile[6][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][14] .is_wysiwyg = "true";
defparam \rfile[6][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N29
dffeas \rfile[4][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][14] .is_wysiwyg = "true";
defparam \rfile[4][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N2
cycloneive_lcell_comb \rfile[5][14]~feeder (
// Equation(s):
// \rfile[5][14]~feeder_combout  = \wdat_WB[14]~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_14),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[5][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[5][14]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[5][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N3
dffeas \rfile[5][14] (
	.clk(!CLK),
	.d(\rfile[5][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][14] .is_wysiwyg = "true";
defparam \rfile[5][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N28
cycloneive_lcell_comb \Mux49~10 (
// Equation(s):
// \Mux49~10_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][14]~q ))) # (!instruction_D[16] & (\rfile[4][14]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][14]~q ),
	.datad(\rfile[5][14]~q ),
	.cin(gnd),
	.combout(\Mux49~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~10 .lut_mask = 16'hDC98;
defparam \Mux49~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N16
cycloneive_lcell_comb \Mux49~11 (
// Equation(s):
// \Mux49~11_combout  = (\Mux49~10_combout  & ((\rfile[7][14]~q ) # ((!instruction_D[17])))) # (!\Mux49~10_combout  & (((\rfile[6][14]~q  & instruction_D[17]))))

	.dataa(\rfile[7][14]~q ),
	.datab(\rfile[6][14]~q ),
	.datac(\Mux49~10_combout ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux49~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~11 .lut_mask = 16'hACF0;
defparam \Mux49~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N21
dffeas \rfile[30][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][13] .is_wysiwyg = "true";
defparam \rfile[30][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y30_N7
dffeas \rfile[22][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][13] .is_wysiwyg = "true";
defparam \rfile[22][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N19
dffeas \rfile[18][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][13] .is_wysiwyg = "true";
defparam \rfile[18][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N25
dffeas \rfile[26][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][13] .is_wysiwyg = "true";
defparam \rfile[26][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N18
cycloneive_lcell_comb \Mux50~2 (
// Equation(s):
// \Mux50~2_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[26][13]~q ))) # (!instruction_D[19] & (\rfile[18][13]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[18][13]~q ),
	.datad(\rfile[26][13]~q ),
	.cin(gnd),
	.combout(\Mux50~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~2 .lut_mask = 16'hDC98;
defparam \Mux50~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N6
cycloneive_lcell_comb \Mux50~3 (
// Equation(s):
// \Mux50~3_combout  = (instruction_D[18] & ((\Mux50~2_combout  & (\rfile[30][13]~q )) # (!\Mux50~2_combout  & ((\rfile[22][13]~q ))))) # (!instruction_D[18] & (((\Mux50~2_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[30][13]~q ),
	.datac(\rfile[22][13]~q ),
	.datad(\Mux50~2_combout ),
	.cin(gnd),
	.combout(\Mux50~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~3 .lut_mask = 16'hDDA0;
defparam \Mux50~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y32_N29
dffeas \rfile[28][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][13] .is_wysiwyg = "true";
defparam \rfile[28][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N5
dffeas \rfile[16][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][13] .is_wysiwyg = "true";
defparam \rfile[16][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N11
dffeas \rfile[24][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][13] .is_wysiwyg = "true";
defparam \rfile[24][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N10
cycloneive_lcell_comb \Mux50~4 (
// Equation(s):
// \Mux50~4_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[24][13]~q ))) # (!instruction_D[19] & (\rfile[16][13]~q ))))

	.dataa(instruction_D_18),
	.datab(\rfile[16][13]~q ),
	.datac(\rfile[24][13]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux50~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~4 .lut_mask = 16'hFA44;
defparam \Mux50~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N28
cycloneive_lcell_comb \Mux50~5 (
// Equation(s):
// \Mux50~5_combout  = (instruction_D[18] & ((\Mux50~4_combout  & ((\rfile[28][13]~q ))) # (!\Mux50~4_combout  & (\rfile[20][13]~q )))) # (!instruction_D[18] & (((\Mux50~4_combout ))))

	.dataa(\rfile[20][13]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[28][13]~q ),
	.datad(\Mux50~4_combout ),
	.cin(gnd),
	.combout(\Mux50~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~5 .lut_mask = 16'hF388;
defparam \Mux50~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N20
cycloneive_lcell_comb \Mux50~6 (
// Equation(s):
// \Mux50~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\Mux50~3_combout )) # (!instruction_D[17] & ((\Mux50~5_combout )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux50~3_combout ),
	.datad(\Mux50~5_combout ),
	.cin(gnd),
	.combout(\Mux50~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~6 .lut_mask = 16'hD9C8;
defparam \Mux50~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N16
cycloneive_lcell_comb \rfile[25][13]~feeder (
// Equation(s):
// \rfile[25][13]~feeder_combout  = \wdat_WB[13]~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_13),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[25][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[25][13]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[25][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N17
dffeas \rfile[25][13] (
	.clk(!CLK),
	.d(\rfile[25][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][13] .is_wysiwyg = "true";
defparam \rfile[25][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N31
dffeas \rfile[29][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][13] .is_wysiwyg = "true";
defparam \rfile[29][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N13
dffeas \rfile[21][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][13] .is_wysiwyg = "true";
defparam \rfile[21][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N25
dffeas \rfile[17][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][13] .is_wysiwyg = "true";
defparam \rfile[17][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N12
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[21][13]~q )) # (!instruction_D[18] & ((\rfile[17][13]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[21][13]~q ),
	.datad(\rfile[17][13]~q ),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'hD9C8;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N30
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (instruction_D[19] & ((\Mux50~0_combout  & ((\rfile[29][13]~q ))) # (!\Mux50~0_combout  & (\rfile[25][13]~q )))) # (!instruction_D[19] & (((\Mux50~0_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[25][13]~q ),
	.datac(\rfile[29][13]~q ),
	.datad(\Mux50~0_combout ),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hF588;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y28_N18
cycloneive_lcell_comb \rfile[27][13]~feeder (
// Equation(s):
// \rfile[27][13]~feeder_combout  = \wdat_WB[13]~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_13),
	.cin(gnd),
	.combout(\rfile[27][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[27][13]~feeder .lut_mask = 16'hFF00;
defparam \rfile[27][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y28_N19
dffeas \rfile[27][13] (
	.clk(!CLK),
	.d(\rfile[27][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][13] .is_wysiwyg = "true";
defparam \rfile[27][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y28_N3
dffeas \rfile[31][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][13] .is_wysiwyg = "true";
defparam \rfile[31][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N1
dffeas \rfile[23][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][13] .is_wysiwyg = "true";
defparam \rfile[23][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N11
dffeas \rfile[19][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][13] .is_wysiwyg = "true";
defparam \rfile[19][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N0
cycloneive_lcell_comb \Mux50~7 (
// Equation(s):
// \Mux50~7_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[23][13]~q )) # (!instruction_D[18] & ((\rfile[19][13]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[23][13]~q ),
	.datad(\rfile[19][13]~q ),
	.cin(gnd),
	.combout(\Mux50~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~7 .lut_mask = 16'hD9C8;
defparam \Mux50~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N2
cycloneive_lcell_comb \Mux50~8 (
// Equation(s):
// \Mux50~8_combout  = (instruction_D[19] & ((\Mux50~7_combout  & ((\rfile[31][13]~q ))) # (!\Mux50~7_combout  & (\rfile[27][13]~q )))) # (!instruction_D[19] & (((\Mux50~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[27][13]~q ),
	.datac(\rfile[31][13]~q ),
	.datad(\Mux50~7_combout ),
	.cin(gnd),
	.combout(\Mux50~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~8 .lut_mask = 16'hF588;
defparam \Mux50~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y30_N17
dffeas \rfile[1][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][13] .is_wysiwyg = "true";
defparam \rfile[1][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N18
cycloneive_lcell_comb \rfile[3][13]~feeder (
// Equation(s):
// \rfile[3][13]~feeder_combout  = \wdat_WB[13]~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_13),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[3][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[3][13]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[3][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y30_N19
dffeas \rfile[3][13] (
	.clk(!CLK),
	.d(\rfile[3][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][13] .is_wysiwyg = "true";
defparam \rfile[3][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N16
cycloneive_lcell_comb \Mux50~14 (
// Equation(s):
// \Mux50~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][13]~q ))) # (!instruction_D[17] & (\rfile[1][13]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[1][13]~q ),
	.datad(\rfile[3][13]~q ),
	.cin(gnd),
	.combout(\Mux50~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~14 .lut_mask = 16'hC840;
defparam \Mux50~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N27
dffeas \rfile[2][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][13] .is_wysiwyg = "true";
defparam \rfile[2][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N26
cycloneive_lcell_comb \Mux50~15 (
// Equation(s):
// \Mux50~15_combout  = (\Mux50~14_combout ) # ((instruction_D[17] & (\rfile[2][13]~q  & !instruction_D[16])))

	.dataa(instruction_D_17),
	.datab(\Mux50~14_combout ),
	.datac(\rfile[2][13]~q ),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux50~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~15 .lut_mask = 16'hCCEC;
defparam \Mux50~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N29
dffeas \rfile[6][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][13] .is_wysiwyg = "true";
defparam \rfile[6][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N17
dffeas \rfile[4][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][13] .is_wysiwyg = "true";
defparam \rfile[4][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N25
dffeas \rfile[5][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][13] .is_wysiwyg = "true";
defparam \rfile[5][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N16
cycloneive_lcell_comb \Mux50~12 (
// Equation(s):
// \Mux50~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][13]~q ))) # (!instruction_D[16] & (\rfile[4][13]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][13]~q ),
	.datad(\rfile[5][13]~q ),
	.cin(gnd),
	.combout(\Mux50~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~12 .lut_mask = 16'hDC98;
defparam \Mux50~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N28
cycloneive_lcell_comb \Mux50~13 (
// Equation(s):
// \Mux50~13_combout  = (instruction_D[17] & ((\Mux50~12_combout  & (\rfile[7][13]~q )) # (!\Mux50~12_combout  & ((\rfile[6][13]~q ))))) # (!instruction_D[17] & (((\Mux50~12_combout ))))

	.dataa(\rfile[7][13]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[6][13]~q ),
	.datad(\Mux50~12_combout ),
	.cin(gnd),
	.combout(\Mux50~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~13 .lut_mask = 16'hBBC0;
defparam \Mux50~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N24
cycloneive_lcell_comb \Mux50~16 (
// Equation(s):
// \Mux50~16_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\Mux50~13_combout )))) # (!instruction_D[18] & (!instruction_D[19] & (\Mux50~15_combout )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\Mux50~15_combout ),
	.datad(\Mux50~13_combout ),
	.cin(gnd),
	.combout(\Mux50~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~16 .lut_mask = 16'hBA98;
defparam \Mux50~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N11
dffeas \rfile[11][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][13] .is_wysiwyg = "true";
defparam \rfile[11][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N25
dffeas \rfile[9][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][13] .is_wysiwyg = "true";
defparam \rfile[9][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N19
dffeas \rfile[8][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][13] .is_wysiwyg = "true";
defparam \rfile[8][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N21
dffeas \rfile[10][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][13] .is_wysiwyg = "true";
defparam \rfile[10][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N18
cycloneive_lcell_comb \Mux50~10 (
// Equation(s):
// \Mux50~10_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][13]~q ))) # (!instruction_D[17] & (\rfile[8][13]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[8][13]~q ),
	.datad(\rfile[10][13]~q ),
	.cin(gnd),
	.combout(\Mux50~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~10 .lut_mask = 16'hDC98;
defparam \Mux50~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N24
cycloneive_lcell_comb \Mux50~11 (
// Equation(s):
// \Mux50~11_combout  = (instruction_D[16] & ((\Mux50~10_combout  & (\rfile[11][13]~q )) # (!\Mux50~10_combout  & ((\rfile[9][13]~q ))))) # (!instruction_D[16] & (((\Mux50~10_combout ))))

	.dataa(\rfile[11][13]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[9][13]~q ),
	.datad(\Mux50~10_combout ),
	.cin(gnd),
	.combout(\Mux50~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~11 .lut_mask = 16'hBBC0;
defparam \Mux50~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N12
cycloneive_lcell_comb \rfile[15][13]~feeder (
// Equation(s):
// \rfile[15][13]~feeder_combout  = \wdat_WB[13]~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_13),
	.cin(gnd),
	.combout(\rfile[15][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][13]~feeder .lut_mask = 16'hFF00;
defparam \rfile[15][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N13
dffeas \rfile[15][13] (
	.clk(!CLK),
	.d(\rfile[15][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][13] .is_wysiwyg = "true";
defparam \rfile[15][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N4
cycloneive_lcell_comb \rfile[14][13]~feeder (
// Equation(s):
// \rfile[14][13]~feeder_combout  = \wdat_WB[13]~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_13),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[14][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][13]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[14][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N5
dffeas \rfile[14][13] (
	.clk(!CLK),
	.d(\rfile[14][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][13] .is_wysiwyg = "true";
defparam \rfile[14][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N19
dffeas \rfile[13][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][13] .is_wysiwyg = "true";
defparam \rfile[13][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N9
dffeas \rfile[12][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][13] .is_wysiwyg = "true";
defparam \rfile[12][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N18
cycloneive_lcell_comb \Mux50~17 (
// Equation(s):
// \Mux50~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][13]~q )))) # (!instruction_D[16] & (!instruction_D[17] & ((\rfile[12][13]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[13][13]~q ),
	.datad(\rfile[12][13]~q ),
	.cin(gnd),
	.combout(\Mux50~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~17 .lut_mask = 16'hB9A8;
defparam \Mux50~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N8
cycloneive_lcell_comb \Mux50~18 (
// Equation(s):
// \Mux50~18_combout  = (instruction_D[17] & ((\Mux50~17_combout  & (\rfile[15][13]~q )) # (!\Mux50~17_combout  & ((\rfile[14][13]~q ))))) # (!instruction_D[17] & (((\Mux50~17_combout ))))

	.dataa(\rfile[15][13]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[14][13]~q ),
	.datad(\Mux50~17_combout ),
	.cin(gnd),
	.combout(\Mux50~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~18 .lut_mask = 16'hBBC0;
defparam \Mux50~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y29_N31
dffeas \rfile[31][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][12] .is_wysiwyg = "true";
defparam \rfile[31][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N5
dffeas \rfile[19][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][12] .is_wysiwyg = "true";
defparam \rfile[19][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N7
dffeas \rfile[27][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][12] .is_wysiwyg = "true";
defparam \rfile[27][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N6
cycloneive_lcell_comb \Mux51~7 (
// Equation(s):
// \Mux51~7_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[27][12]~q ))) # (!instruction_D[19] & (\rfile[19][12]~q ))))

	.dataa(instruction_D_18),
	.datab(\rfile[19][12]~q ),
	.datac(\rfile[27][12]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux51~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~7 .lut_mask = 16'hFA44;
defparam \Mux51~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y29_N1
dffeas \rfile[23][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][12] .is_wysiwyg = "true";
defparam \rfile[23][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N0
cycloneive_lcell_comb \Mux51~8 (
// Equation(s):
// \Mux51~8_combout  = (\Mux51~7_combout  & ((\rfile[31][12]~q ) # ((!instruction_D[18])))) # (!\Mux51~7_combout  & (((\rfile[23][12]~q  & instruction_D[18]))))

	.dataa(\rfile[31][12]~q ),
	.datab(\Mux51~7_combout ),
	.datac(\rfile[23][12]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux51~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~8 .lut_mask = 16'hB8CC;
defparam \Mux51~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N26
cycloneive_lcell_comb \rfile[21][12]~feeder (
// Equation(s):
// \rfile[21][12]~feeder_combout  = \wdat_WB[12]~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[21][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][12]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[21][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N27
dffeas \rfile[21][12] (
	.clk(!CLK),
	.d(\rfile[21][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][12] .is_wysiwyg = "true";
defparam \rfile[21][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N9
dffeas \rfile[29][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][12] .is_wysiwyg = "true";
defparam \rfile[29][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y30_N15
dffeas \rfile[17][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][12] .is_wysiwyg = "true";
defparam \rfile[17][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y30_N21
dffeas \rfile[25][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][12] .is_wysiwyg = "true";
defparam \rfile[25][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N14
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[25][12]~q ))) # (!instruction_D[19] & (\rfile[17][12]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[17][12]~q ),
	.datad(\rfile[25][12]~q ),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'hDC98;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N8
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (instruction_D[18] & ((\Mux51~0_combout  & ((\rfile[29][12]~q ))) # (!\Mux51~0_combout  & (\rfile[21][12]~q )))) # (!instruction_D[18] & (((\Mux51~0_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[21][12]~q ),
	.datac(\rfile[29][12]~q ),
	.datad(\Mux51~0_combout ),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hF588;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y30_N17
dffeas \rfile[28][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][12] .is_wysiwyg = "true";
defparam \rfile[28][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N22
cycloneive_lcell_comb \rfile[20][12]~feeder (
// Equation(s):
// \rfile[20][12]~feeder_combout  = \wdat_WB[12]~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_12),
	.cin(gnd),
	.combout(\rfile[20][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[20][12]~feeder .lut_mask = 16'hFF00;
defparam \rfile[20][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y30_N23
dffeas \rfile[20][12] (
	.clk(!CLK),
	.d(\rfile[20][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][12] .is_wysiwyg = "true";
defparam \rfile[20][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N24
cycloneive_lcell_comb \rfile[16][12]~feeder (
// Equation(s):
// \rfile[16][12]~feeder_combout  = \wdat_WB[12]~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_12),
	.cin(gnd),
	.combout(\rfile[16][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[16][12]~feeder .lut_mask = 16'hFF00;
defparam \rfile[16][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y30_N25
dffeas \rfile[16][12] (
	.clk(!CLK),
	.d(\rfile[16][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][12] .is_wysiwyg = "true";
defparam \rfile[16][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N6
cycloneive_lcell_comb \Mux51~4 (
// Equation(s):
// \Mux51~4_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[20][12]~q )) # (!instruction_D[18] & ((\rfile[16][12]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[20][12]~q ),
	.datad(\rfile[16][12]~q ),
	.cin(gnd),
	.combout(\Mux51~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~4 .lut_mask = 16'hD9C8;
defparam \Mux51~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N16
cycloneive_lcell_comb \Mux51~5 (
// Equation(s):
// \Mux51~5_combout  = (instruction_D[19] & ((\Mux51~4_combout  & ((\rfile[28][12]~q ))) # (!\Mux51~4_combout  & (\rfile[24][12]~q )))) # (!instruction_D[19] & (((\Mux51~4_combout ))))

	.dataa(\rfile[24][12]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[28][12]~q ),
	.datad(\Mux51~4_combout ),
	.cin(gnd),
	.combout(\Mux51~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~5 .lut_mask = 16'hF388;
defparam \Mux51~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y36_N5
dffeas \rfile[26][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][12] .is_wysiwyg = "true";
defparam \rfile[26][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y34_N19
dffeas \rfile[22][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][12] .is_wysiwyg = "true";
defparam \rfile[22][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y34_N1
dffeas \rfile[18][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][12] .is_wysiwyg = "true";
defparam \rfile[18][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N18
cycloneive_lcell_comb \Mux51~2 (
// Equation(s):
// \Mux51~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[22][12]~q )) # (!instruction_D[18] & ((\rfile[18][12]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[22][12]~q ),
	.datad(\rfile[18][12]~q ),
	.cin(gnd),
	.combout(\Mux51~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~2 .lut_mask = 16'hD9C8;
defparam \Mux51~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N4
cycloneive_lcell_comb \Mux51~3 (
// Equation(s):
// \Mux51~3_combout  = (instruction_D[19] & ((\Mux51~2_combout  & (\rfile[30][12]~q )) # (!\Mux51~2_combout  & ((\rfile[26][12]~q ))))) # (!instruction_D[19] & (((\Mux51~2_combout ))))

	.dataa(\rfile[30][12]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[26][12]~q ),
	.datad(\Mux51~2_combout ),
	.cin(gnd),
	.combout(\Mux51~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~3 .lut_mask = 16'hBBC0;
defparam \Mux51~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N2
cycloneive_lcell_comb \Mux51~6 (
// Equation(s):
// \Mux51~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\Mux51~3_combout ))) # (!instruction_D[17] & (\Mux51~5_combout ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux51~5_combout ),
	.datad(\Mux51~3_combout ),
	.cin(gnd),
	.combout(\Mux51~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~6 .lut_mask = 16'hDC98;
defparam \Mux51~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N22
cycloneive_lcell_comb \rfile[15][12]~feeder (
// Equation(s):
// \rfile[15][12]~feeder_combout  = \wdat_WB[12]~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_12),
	.cin(gnd),
	.combout(\rfile[15][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][12]~feeder .lut_mask = 16'hFF00;
defparam \rfile[15][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N23
dffeas \rfile[15][12] (
	.clk(!CLK),
	.d(\rfile[15][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][12] .is_wysiwyg = "true";
defparam \rfile[15][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N23
dffeas \rfile[14][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][12] .is_wysiwyg = "true";
defparam \rfile[14][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N17
dffeas \rfile[13][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][12] .is_wysiwyg = "true";
defparam \rfile[13][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N23
dffeas \rfile[12][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][12] .is_wysiwyg = "true";
defparam \rfile[12][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N16
cycloneive_lcell_comb \Mux51~17 (
// Equation(s):
// \Mux51~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][12]~q )))) # (!instruction_D[16] & (!instruction_D[17] & ((\rfile[12][12]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[13][12]~q ),
	.datad(\rfile[12][12]~q ),
	.cin(gnd),
	.combout(\Mux51~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~17 .lut_mask = 16'hB9A8;
defparam \Mux51~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N22
cycloneive_lcell_comb \Mux51~18 (
// Equation(s):
// \Mux51~18_combout  = (instruction_D[17] & ((\Mux51~17_combout  & (\rfile[15][12]~q )) # (!\Mux51~17_combout  & ((\rfile[14][12]~q ))))) # (!instruction_D[17] & (((\Mux51~17_combout ))))

	.dataa(\rfile[15][12]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[14][12]~q ),
	.datad(\Mux51~17_combout ),
	.cin(gnd),
	.combout(\Mux51~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~18 .lut_mask = 16'hBBC0;
defparam \Mux51~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N13
dffeas \rfile[5][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][12] .is_wysiwyg = "true";
defparam \rfile[5][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N12
cycloneive_lcell_comb \Mux51~10 (
// Equation(s):
// \Mux51~10_combout  = (instruction_D[16] & (((\rfile[5][12]~q ) # (instruction_D[17])))) # (!instruction_D[16] & (\rfile[4][12]~q  & ((!instruction_D[17]))))

	.dataa(\rfile[4][12]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[5][12]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux51~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~10 .lut_mask = 16'hCCE2;
defparam \Mux51~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N27
dffeas \rfile[6][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][12] .is_wysiwyg = "true";
defparam \rfile[6][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N21
dffeas \rfile[7][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][12] .is_wysiwyg = "true";
defparam \rfile[7][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N26
cycloneive_lcell_comb \Mux51~11 (
// Equation(s):
// \Mux51~11_combout  = (\Mux51~10_combout  & (((\rfile[7][12]~q )) # (!instruction_D[17]))) # (!\Mux51~10_combout  & (instruction_D[17] & (\rfile[6][12]~q )))

	.dataa(\Mux51~10_combout ),
	.datab(instruction_D_17),
	.datac(\rfile[6][12]~q ),
	.datad(\rfile[7][12]~q ),
	.cin(gnd),
	.combout(\Mux51~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~11 .lut_mask = 16'hEA62;
defparam \Mux51~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N27
dffeas \rfile[2][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][12] .is_wysiwyg = "true";
defparam \rfile[2][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N29
dffeas \rfile[3][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][12] .is_wysiwyg = "true";
defparam \rfile[3][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N3
dffeas \rfile[1][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][12] .is_wysiwyg = "true";
defparam \rfile[1][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N28
cycloneive_lcell_comb \Mux51~14 (
// Equation(s):
// \Mux51~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][12]~q )) # (!instruction_D[17] & ((\rfile[1][12]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[3][12]~q ),
	.datad(\rfile[1][12]~q ),
	.cin(gnd),
	.combout(\Mux51~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~14 .lut_mask = 16'hA280;
defparam \Mux51~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N26
cycloneive_lcell_comb \Mux51~15 (
// Equation(s):
// \Mux51~15_combout  = (\Mux51~14_combout ) # ((instruction_D[17] & (!instruction_D[16] & \rfile[2][12]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[2][12]~q ),
	.datad(\Mux51~14_combout ),
	.cin(gnd),
	.combout(\Mux51~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~15 .lut_mask = 16'hFF20;
defparam \Mux51~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N23
dffeas \rfile[11][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][12] .is_wysiwyg = "true";
defparam \rfile[11][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N24
cycloneive_lcell_comb \rfile[9][12]~feeder (
// Equation(s):
// \rfile[9][12]~feeder_combout  = \wdat_WB[12]~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_12),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[9][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][12]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[9][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N25
dffeas \rfile[9][12] (
	.clk(!CLK),
	.d(\rfile[9][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][12] .is_wysiwyg = "true";
defparam \rfile[9][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N22
cycloneive_lcell_comb \Mux51~13 (
// Equation(s):
// \Mux51~13_combout  = (\Mux51~12_combout  & (((\rfile[11][12]~q )) # (!instruction_D[16]))) # (!\Mux51~12_combout  & (instruction_D[16] & ((\rfile[9][12]~q ))))

	.dataa(\Mux51~12_combout ),
	.datab(instruction_D_16),
	.datac(\rfile[11][12]~q ),
	.datad(\rfile[9][12]~q ),
	.cin(gnd),
	.combout(\Mux51~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~13 .lut_mask = 16'hE6A2;
defparam \Mux51~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N28
cycloneive_lcell_comb \Mux51~16 (
// Equation(s):
// \Mux51~16_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\Mux51~13_combout ))) # (!instruction_D[19] & (\Mux51~15_combout ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\Mux51~15_combout ),
	.datad(\Mux51~13_combout ),
	.cin(gnd),
	.combout(\Mux51~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~16 .lut_mask = 16'hDC98;
defparam \Mux51~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N3
dffeas \rfile[17][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][9] .is_wysiwyg = "true";
defparam \rfile[17][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y30_N5
dffeas \rfile[21][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][9] .is_wysiwyg = "true";
defparam \rfile[21][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N2
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[21][9]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[17][9]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[17][9]~q ),
	.datad(\rfile[21][9]~q ),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'hBA98;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N21
dffeas \rfile[29][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][9] .is_wysiwyg = "true";
defparam \rfile[29][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N7
dffeas \rfile[25][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][9] .is_wysiwyg = "true";
defparam \rfile[25][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N20
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (instruction_D[19] & ((\Mux54~0_combout  & (\rfile[29][9]~q )) # (!\Mux54~0_combout  & ((\rfile[25][9]~q ))))) # (!instruction_D[19] & (\Mux54~0_combout ))

	.dataa(instruction_D_19),
	.datab(\Mux54~0_combout ),
	.datac(\rfile[29][9]~q ),
	.datad(\rfile[25][9]~q ),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hE6C4;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y27_N0
cycloneive_lcell_comb \rfile[27][9]~feeder (
// Equation(s):
// \rfile[27][9]~feeder_combout  = \wdat_WB[9]~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_9),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[27][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[27][9]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[27][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y27_N1
dffeas \rfile[27][9] (
	.clk(!CLK),
	.d(\rfile[27][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][9] .is_wysiwyg = "true";
defparam \rfile[27][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y28_N27
dffeas \rfile[31][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][9] .is_wysiwyg = "true";
defparam \rfile[31][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N28
cycloneive_lcell_comb \rfile[23][9]~feeder (
// Equation(s):
// \rfile[23][9]~feeder_combout  = \wdat_WB[9]~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_9),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[23][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[23][9]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[23][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y31_N29
dffeas \rfile[23][9] (
	.clk(!CLK),
	.d(\rfile[23][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][9] .is_wysiwyg = "true";
defparam \rfile[23][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y28_N29
dffeas \rfile[19][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][9] .is_wysiwyg = "true";
defparam \rfile[19][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N28
cycloneive_lcell_comb \Mux54~7 (
// Equation(s):
// \Mux54~7_combout  = (instruction_D[19] & (((instruction_D[18])))) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[23][9]~q )) # (!instruction_D[18] & ((\rfile[19][9]~q )))))

	.dataa(instruction_D_19),
	.datab(\rfile[23][9]~q ),
	.datac(\rfile[19][9]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux54~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~7 .lut_mask = 16'hEE50;
defparam \Mux54~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N20
cycloneive_lcell_comb \Mux54~8 (
// Equation(s):
// \Mux54~8_combout  = (instruction_D[19] & ((\Mux54~7_combout  & ((\rfile[31][9]~q ))) # (!\Mux54~7_combout  & (\rfile[27][9]~q )))) # (!instruction_D[19] & (((\Mux54~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[27][9]~q ),
	.datac(\rfile[31][9]~q ),
	.datad(\Mux54~7_combout ),
	.cin(gnd),
	.combout(\Mux54~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~8 .lut_mask = 16'hF588;
defparam \Mux54~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N5
dffeas \rfile[30][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][9] .is_wysiwyg = "true";
defparam \rfile[30][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y34_N7
dffeas \rfile[22][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][9] .is_wysiwyg = "true";
defparam \rfile[22][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y36_N29
dffeas \rfile[26][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][9] .is_wysiwyg = "true";
defparam \rfile[26][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y36_N29
dffeas \rfile[18][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][9] .is_wysiwyg = "true";
defparam \rfile[18][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N28
cycloneive_lcell_comb \Mux54~2 (
// Equation(s):
// \Mux54~2_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[26][9]~q )) # (!instruction_D[19] & ((\rfile[18][9]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[26][9]~q ),
	.datad(\rfile[18][9]~q ),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~2 .lut_mask = 16'hD9C8;
defparam \Mux54~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N6
cycloneive_lcell_comb \Mux54~3 (
// Equation(s):
// \Mux54~3_combout  = (instruction_D[18] & ((\Mux54~2_combout  & (\rfile[30][9]~q )) # (!\Mux54~2_combout  & ((\rfile[22][9]~q ))))) # (!instruction_D[18] & (((\Mux54~2_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[30][9]~q ),
	.datac(\rfile[22][9]~q ),
	.datad(\Mux54~2_combout ),
	.cin(gnd),
	.combout(\Mux54~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~3 .lut_mask = 16'hDDA0;
defparam \Mux54~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y32_N15
dffeas \rfile[28][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][9] .is_wysiwyg = "true";
defparam \rfile[28][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N25
dffeas \rfile[16][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][9] .is_wysiwyg = "true";
defparam \rfile[16][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N7
dffeas \rfile[24][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][9] .is_wysiwyg = "true";
defparam \rfile[24][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N24
cycloneive_lcell_comb \Mux54~4 (
// Equation(s):
// \Mux54~4_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[24][9]~q ))) # (!instruction_D[19] & (\rfile[16][9]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[16][9]~q ),
	.datad(\rfile[24][9]~q ),
	.cin(gnd),
	.combout(\Mux54~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~4 .lut_mask = 16'hDC98;
defparam \Mux54~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N14
cycloneive_lcell_comb \Mux54~5 (
// Equation(s):
// \Mux54~5_combout  = (instruction_D[18] & ((\Mux54~4_combout  & ((\rfile[28][9]~q ))) # (!\Mux54~4_combout  & (\rfile[20][9]~q )))) # (!instruction_D[18] & (((\Mux54~4_combout ))))

	.dataa(\rfile[20][9]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[28][9]~q ),
	.datad(\Mux54~4_combout ),
	.cin(gnd),
	.combout(\Mux54~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~5 .lut_mask = 16'hF388;
defparam \Mux54~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N6
cycloneive_lcell_comb \Mux54~6 (
// Equation(s):
// \Mux54~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\Mux54~3_combout )) # (!instruction_D[17] & ((\Mux54~5_combout )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux54~3_combout ),
	.datad(\Mux54~5_combout ),
	.cin(gnd),
	.combout(\Mux54~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~6 .lut_mask = 16'hD9C8;
defparam \Mux54~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N8
cycloneive_lcell_comb \rfile[15][9]~feeder (
// Equation(s):
// \rfile[15][9]~feeder_combout  = \wdat_WB[9]~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_9),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[15][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][9]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[15][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N9
dffeas \rfile[15][9] (
	.clk(!CLK),
	.d(\rfile[15][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][9] .is_wysiwyg = "true";
defparam \rfile[15][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N28
cycloneive_lcell_comb \rfile[14][9]~feeder (
// Equation(s):
// \rfile[14][9]~feeder_combout  = \wdat_WB[9]~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_9),
	.cin(gnd),
	.combout(\rfile[14][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][9]~feeder .lut_mask = 16'hFF00;
defparam \rfile[14][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N29
dffeas \rfile[14][9] (
	.clk(!CLK),
	.d(\rfile[14][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][9] .is_wysiwyg = "true";
defparam \rfile[14][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N7
dffeas \rfile[12][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][9] .is_wysiwyg = "true";
defparam \rfile[12][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N9
dffeas \rfile[13][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][9] .is_wysiwyg = "true";
defparam \rfile[13][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N6
cycloneive_lcell_comb \Mux54~17 (
// Equation(s):
// \Mux54~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][9]~q ))) # (!instruction_D[16] & (\rfile[12][9]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][9]~q ),
	.datad(\rfile[13][9]~q ),
	.cin(gnd),
	.combout(\Mux54~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~17 .lut_mask = 16'hDC98;
defparam \Mux54~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N30
cycloneive_lcell_comb \Mux54~18 (
// Equation(s):
// \Mux54~18_combout  = (instruction_D[17] & ((\Mux54~17_combout  & (\rfile[15][9]~q )) # (!\Mux54~17_combout  & ((\rfile[14][9]~q ))))) # (!instruction_D[17] & (((\Mux54~17_combout ))))

	.dataa(\rfile[15][9]~q ),
	.datab(\rfile[14][9]~q ),
	.datac(instruction_D_17),
	.datad(\Mux54~17_combout ),
	.cin(gnd),
	.combout(\Mux54~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~18 .lut_mask = 16'hAFC0;
defparam \Mux54~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N31
dffeas \rfile[11][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][9] .is_wysiwyg = "true";
defparam \rfile[11][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N29
dffeas \rfile[9][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][9] .is_wysiwyg = "true";
defparam \rfile[9][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N3
dffeas \rfile[8][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][9] .is_wysiwyg = "true";
defparam \rfile[8][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N13
dffeas \rfile[10][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][9] .is_wysiwyg = "true";
defparam \rfile[10][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N2
cycloneive_lcell_comb \Mux54~10 (
// Equation(s):
// \Mux54~10_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][9]~q ))) # (!instruction_D[17] & (\rfile[8][9]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[8][9]~q ),
	.datad(\rfile[10][9]~q ),
	.cin(gnd),
	.combout(\Mux54~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~10 .lut_mask = 16'hDC98;
defparam \Mux54~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N28
cycloneive_lcell_comb \Mux54~11 (
// Equation(s):
// \Mux54~11_combout  = (instruction_D[16] & ((\Mux54~10_combout  & (\rfile[11][9]~q )) # (!\Mux54~10_combout  & ((\rfile[9][9]~q ))))) # (!instruction_D[16] & (((\Mux54~10_combout ))))

	.dataa(\rfile[11][9]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[9][9]~q ),
	.datad(\Mux54~10_combout ),
	.cin(gnd),
	.combout(\Mux54~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~11 .lut_mask = 16'hBBC0;
defparam \Mux54~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y27_N19
dffeas \rfile[1][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][9] .is_wysiwyg = "true";
defparam \rfile[1][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N25
dffeas \rfile[3][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][9] .is_wysiwyg = "true";
defparam \rfile[3][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N18
cycloneive_lcell_comb \Mux54~14 (
// Equation(s):
// \Mux54~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][9]~q ))) # (!instruction_D[17] & (\rfile[1][9]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[1][9]~q ),
	.datad(\rfile[3][9]~q ),
	.cin(gnd),
	.combout(\Mux54~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~14 .lut_mask = 16'hA820;
defparam \Mux54~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N26
cycloneive_lcell_comb \Mux54~15 (
// Equation(s):
// \Mux54~15_combout  = (\Mux54~14_combout ) # ((\rfile[2][9]~q  & (instruction_D[17] & !instruction_D[16])))

	.dataa(\rfile[2][9]~q ),
	.datab(instruction_D_17),
	.datac(instruction_D_16),
	.datad(\Mux54~14_combout ),
	.cin(gnd),
	.combout(\Mux54~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~15 .lut_mask = 16'hFF08;
defparam \Mux54~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N19
dffeas \rfile[6][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][9] .is_wysiwyg = "true";
defparam \rfile[6][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y28_N31
dffeas \rfile[7][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][9] .is_wysiwyg = "true";
defparam \rfile[7][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N18
cycloneive_lcell_comb \Mux54~13 (
// Equation(s):
// \Mux54~13_combout  = (\Mux54~12_combout  & (((\rfile[7][9]~q )) # (!instruction_D[17]))) # (!\Mux54~12_combout  & (instruction_D[17] & (\rfile[6][9]~q )))

	.dataa(\Mux54~12_combout ),
	.datab(instruction_D_17),
	.datac(\rfile[6][9]~q ),
	.datad(\rfile[7][9]~q ),
	.cin(gnd),
	.combout(\Mux54~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~13 .lut_mask = 16'hEA62;
defparam \Mux54~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N28
cycloneive_lcell_comb \Mux54~16 (
// Equation(s):
// \Mux54~16_combout  = (instruction_D[19] & (((instruction_D[18])))) # (!instruction_D[19] & ((instruction_D[18] & ((\Mux54~13_combout ))) # (!instruction_D[18] & (\Mux54~15_combout ))))

	.dataa(\Mux54~15_combout ),
	.datab(instruction_D_19),
	.datac(instruction_D_18),
	.datad(\Mux54~13_combout ),
	.cin(gnd),
	.combout(\Mux54~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~16 .lut_mask = 16'hF2C2;
defparam \Mux54~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y29_N23
dffeas \rfile[31][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][8] .is_wysiwyg = "true";
defparam \rfile[31][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y29_N5
dffeas \rfile[23][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][8] .is_wysiwyg = "true";
defparam \rfile[23][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N25
dffeas \rfile[19][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][8] .is_wysiwyg = "true";
defparam \rfile[19][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N19
dffeas \rfile[27][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][8] .is_wysiwyg = "true";
defparam \rfile[27][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N24
cycloneive_lcell_comb \Mux55~7 (
// Equation(s):
// \Mux55~7_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[27][8]~q )))) # (!instruction_D[19] & (!instruction_D[18] & (\rfile[19][8]~q )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[19][8]~q ),
	.datad(\rfile[27][8]~q ),
	.cin(gnd),
	.combout(\Mux55~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~7 .lut_mask = 16'hBA98;
defparam \Mux55~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N4
cycloneive_lcell_comb \Mux55~8 (
// Equation(s):
// \Mux55~8_combout  = (instruction_D[18] & ((\Mux55~7_combout  & (\rfile[31][8]~q )) # (!\Mux55~7_combout  & ((\rfile[23][8]~q ))))) # (!instruction_D[18] & (((\Mux55~7_combout ))))

	.dataa(\rfile[31][8]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[23][8]~q ),
	.datad(\Mux55~7_combout ),
	.cin(gnd),
	.combout(\Mux55~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~8 .lut_mask = 16'hBBC0;
defparam \Mux55~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y36_N1
dffeas \rfile[26][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][8] .is_wysiwyg = "true";
defparam \rfile[26][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y35_N1
dffeas \rfile[18][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][8] .is_wysiwyg = "true";
defparam \rfile[18][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y35_N19
dffeas \rfile[22][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][8] .is_wysiwyg = "true";
defparam \rfile[22][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N0
cycloneive_lcell_comb \Mux55~2 (
// Equation(s):
// \Mux55~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[22][8]~q ))) # (!instruction_D[18] & (\rfile[18][8]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][8]~q ),
	.datad(\rfile[22][8]~q ),
	.cin(gnd),
	.combout(\Mux55~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~2 .lut_mask = 16'hDC98;
defparam \Mux55~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N0
cycloneive_lcell_comb \Mux55~3 (
// Equation(s):
// \Mux55~3_combout  = (instruction_D[19] & ((\Mux55~2_combout  & (\rfile[30][8]~q )) # (!\Mux55~2_combout  & ((\rfile[26][8]~q ))))) # (!instruction_D[19] & (((\Mux55~2_combout ))))

	.dataa(\rfile[30][8]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[26][8]~q ),
	.datad(\Mux55~2_combout ),
	.cin(gnd),
	.combout(\Mux55~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~3 .lut_mask = 16'hBBC0;
defparam \Mux55~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y30_N19
dffeas \rfile[24][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][8] .is_wysiwyg = "true";
defparam \rfile[24][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X77_Y30_N22
cycloneive_lcell_comb \rfile[16][8]~feeder (
// Equation(s):
// \rfile[16][8]~feeder_combout  = \wdat_WB[8]~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_8),
	.cin(gnd),
	.combout(\rfile[16][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[16][8]~feeder .lut_mask = 16'hFF00;
defparam \rfile[16][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X77_Y30_N23
dffeas \rfile[16][8] (
	.clk(!CLK),
	.d(\rfile[16][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][8] .is_wysiwyg = "true";
defparam \rfile[16][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X77_Y30_N0
cycloneive_lcell_comb \rfile[20][8]~feeder (
// Equation(s):
// \rfile[20][8]~feeder_combout  = \wdat_WB[8]~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_8),
	.cin(gnd),
	.combout(\rfile[20][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[20][8]~feeder .lut_mask = 16'hFF00;
defparam \rfile[20][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X77_Y30_N1
dffeas \rfile[20][8] (
	.clk(!CLK),
	.d(\rfile[20][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][8] .is_wysiwyg = "true";
defparam \rfile[20][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X77_Y30_N12
cycloneive_lcell_comb \Mux55~4 (
// Equation(s):
// \Mux55~4_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[20][8]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[16][8]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[16][8]~q ),
	.datad(\rfile[20][8]~q ),
	.cin(gnd),
	.combout(\Mux55~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~4 .lut_mask = 16'hBA98;
defparam \Mux55~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N18
cycloneive_lcell_comb \Mux55~5 (
// Equation(s):
// \Mux55~5_combout  = (instruction_D[19] & ((\Mux55~4_combout  & (\rfile[28][8]~q )) # (!\Mux55~4_combout  & ((\rfile[24][8]~q ))))) # (!instruction_D[19] & (((\Mux55~4_combout ))))

	.dataa(\rfile[28][8]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[24][8]~q ),
	.datad(\Mux55~4_combout ),
	.cin(gnd),
	.combout(\Mux55~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~5 .lut_mask = 16'hBBC0;
defparam \Mux55~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N8
cycloneive_lcell_comb \Mux55~6 (
// Equation(s):
// \Mux55~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\Mux55~3_combout )) # (!instruction_D[17] & ((\Mux55~5_combout )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux55~3_combout ),
	.datad(\Mux55~5_combout ),
	.cin(gnd),
	.combout(\Mux55~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~6 .lut_mask = 16'hD9C8;
defparam \Mux55~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N27
dffeas \rfile[29][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][8] .is_wysiwyg = "true";
defparam \rfile[29][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N24
cycloneive_lcell_comb \rfile[21][8]~feeder (
// Equation(s):
// \rfile[21][8]~feeder_combout  = \wdat_WB[8]~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[21][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][8]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[21][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N25
dffeas \rfile[21][8] (
	.clk(!CLK),
	.d(\rfile[21][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][8] .is_wysiwyg = "true";
defparam \rfile[21][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N23
dffeas \rfile[25][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][8] .is_wysiwyg = "true";
defparam \rfile[25][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N7
dffeas \rfile[17][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][8] .is_wysiwyg = "true";
defparam \rfile[17][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N22
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[25][8]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[17][8]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[25][8]~q ),
	.datad(\rfile[17][8]~q ),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'hB9A8;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N2
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (instruction_D[18] & ((\Mux55~0_combout  & (\rfile[29][8]~q )) # (!\Mux55~0_combout  & ((\rfile[21][8]~q ))))) # (!instruction_D[18] & (((\Mux55~0_combout ))))

	.dataa(\rfile[29][8]~q ),
	.datab(\rfile[21][8]~q ),
	.datac(instruction_D_18),
	.datad(\Mux55~0_combout ),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hAFC0;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N27
dffeas \rfile[15][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][8] .is_wysiwyg = "true";
defparam \rfile[15][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N18
cycloneive_lcell_comb \rfile[14][8]~feeder (
// Equation(s):
// \rfile[14][8]~feeder_combout  = \wdat_WB[8]~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[14][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][8]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[14][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N19
dffeas \rfile[14][8] (
	.clk(!CLK),
	.d(\rfile[14][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][8] .is_wysiwyg = "true";
defparam \rfile[14][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N21
dffeas \rfile[12][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][8] .is_wysiwyg = "true";
defparam \rfile[12][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N27
dffeas \rfile[13][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][8] .is_wysiwyg = "true";
defparam \rfile[13][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N20
cycloneive_lcell_comb \Mux55~17 (
// Equation(s):
// \Mux55~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][8]~q ))) # (!instruction_D[16] & (\rfile[12][8]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][8]~q ),
	.datad(\rfile[13][8]~q ),
	.cin(gnd),
	.combout(\Mux55~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~17 .lut_mask = 16'hDC98;
defparam \Mux55~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N4
cycloneive_lcell_comb \Mux55~18 (
// Equation(s):
// \Mux55~18_combout  = (instruction_D[17] & ((\Mux55~17_combout  & (\rfile[15][8]~q )) # (!\Mux55~17_combout  & ((\rfile[14][8]~q ))))) # (!instruction_D[17] & (((\Mux55~17_combout ))))

	.dataa(\rfile[15][8]~q ),
	.datab(\rfile[14][8]~q ),
	.datac(instruction_D_17),
	.datad(\Mux55~17_combout ),
	.cin(gnd),
	.combout(\Mux55~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~18 .lut_mask = 16'hAFC0;
defparam \Mux55~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N2
cycloneive_lcell_comb \rfile[6][8]~feeder (
// Equation(s):
// \rfile[6][8]~feeder_combout  = \wdat_WB[8]~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[6][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][8]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[6][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N3
dffeas \rfile[6][8] (
	.clk(!CLK),
	.d(\rfile[6][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][8] .is_wysiwyg = "true";
defparam \rfile[6][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N5
dffeas \rfile[5][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][8] .is_wysiwyg = "true";
defparam \rfile[5][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N23
dffeas \rfile[4][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][8] .is_wysiwyg = "true";
defparam \rfile[4][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N22
cycloneive_lcell_comb \Mux55~10 (
// Equation(s):
// \Mux55~10_combout  = (instruction_D[17] & (((instruction_D[16])))) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[5][8]~q )) # (!instruction_D[16] & ((\rfile[4][8]~q )))))

	.dataa(instruction_D_17),
	.datab(\rfile[5][8]~q ),
	.datac(\rfile[4][8]~q ),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux55~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~10 .lut_mask = 16'hEE50;
defparam \Mux55~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N0
cycloneive_lcell_comb \rfile[7][8]~feeder (
// Equation(s):
// \rfile[7][8]~feeder_combout  = \wdat_WB[8]~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[7][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[7][8]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[7][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N1
dffeas \rfile[7][8] (
	.clk(!CLK),
	.d(\rfile[7][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][8] .is_wysiwyg = "true";
defparam \rfile[7][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N0
cycloneive_lcell_comb \Mux55~11 (
// Equation(s):
// \Mux55~11_combout  = (instruction_D[17] & ((\Mux55~10_combout  & ((\rfile[7][8]~q ))) # (!\Mux55~10_combout  & (\rfile[6][8]~q )))) # (!instruction_D[17] & (((\Mux55~10_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[6][8]~q ),
	.datac(\Mux55~10_combout ),
	.datad(\rfile[7][8]~q ),
	.cin(gnd),
	.combout(\Mux55~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~11 .lut_mask = 16'hF858;
defparam \Mux55~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N29
dffeas \rfile[11][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][8] .is_wysiwyg = "true";
defparam \rfile[11][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y35_N3
dffeas \rfile[9][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][8] .is_wysiwyg = "true";
defparam \rfile[9][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N15
dffeas \rfile[8][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][8] .is_wysiwyg = "true";
defparam \rfile[8][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N9
dffeas \rfile[10][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][8] .is_wysiwyg = "true";
defparam \rfile[10][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N14
cycloneive_lcell_comb \Mux55~12 (
// Equation(s):
// \Mux55~12_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][8]~q )))) # (!instruction_D[17] & (!instruction_D[16] & (\rfile[8][8]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[8][8]~q ),
	.datad(\rfile[10][8]~q ),
	.cin(gnd),
	.combout(\Mux55~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~12 .lut_mask = 16'hBA98;
defparam \Mux55~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N2
cycloneive_lcell_comb \Mux55~13 (
// Equation(s):
// \Mux55~13_combout  = (instruction_D[16] & ((\Mux55~12_combout  & (\rfile[11][8]~q )) # (!\Mux55~12_combout  & ((\rfile[9][8]~q ))))) # (!instruction_D[16] & (((\Mux55~12_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][8]~q ),
	.datac(\rfile[9][8]~q ),
	.datad(\Mux55~12_combout ),
	.cin(gnd),
	.combout(\Mux55~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~13 .lut_mask = 16'hDDA0;
defparam \Mux55~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N8
cycloneive_lcell_comb \rfile[2][8]~feeder (
// Equation(s):
// \rfile[2][8]~feeder_combout  = \wdat_WB[8]~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[2][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][8]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[2][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N9
dffeas \rfile[2][8] (
	.clk(!CLK),
	.d(\rfile[2][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][8] .is_wysiwyg = "true";
defparam \rfile[2][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N1
dffeas \rfile[3][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][8] .is_wysiwyg = "true";
defparam \rfile[3][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N11
dffeas \rfile[1][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][8] .is_wysiwyg = "true";
defparam \rfile[1][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N0
cycloneive_lcell_comb \Mux55~14 (
// Equation(s):
// \Mux55~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][8]~q )) # (!instruction_D[17] & ((\rfile[1][8]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[3][8]~q ),
	.datad(\rfile[1][8]~q ),
	.cin(gnd),
	.combout(\Mux55~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~14 .lut_mask = 16'hA280;
defparam \Mux55~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N10
cycloneive_lcell_comb \Mux55~15 (
// Equation(s):
// \Mux55~15_combout  = (\Mux55~14_combout ) # ((!instruction_D[16] & (\rfile[2][8]~q  & instruction_D[17])))

	.dataa(instruction_D_16),
	.datab(\rfile[2][8]~q ),
	.datac(instruction_D_17),
	.datad(\Mux55~14_combout ),
	.cin(gnd),
	.combout(\Mux55~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~15 .lut_mask = 16'hFF40;
defparam \Mux55~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N28
cycloneive_lcell_comb \Mux55~16 (
// Equation(s):
// \Mux55~16_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & (\Mux55~13_combout )) # (!instruction_D[19] & ((\Mux55~15_combout )))))

	.dataa(instruction_D_18),
	.datab(\Mux55~13_combout ),
	.datac(\Mux55~15_combout ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux55~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~16 .lut_mask = 16'hEE50;
defparam \Mux55~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y28_N24
cycloneive_lcell_comb \rfile[27][11]~feeder (
// Equation(s):
// \rfile[27][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[27][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[27][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[27][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y28_N25
dffeas \rfile[27][11] (
	.clk(!CLK),
	.d(\rfile[27][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][11] .is_wysiwyg = "true";
defparam \rfile[27][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y28_N7
dffeas \rfile[31][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][11] .is_wysiwyg = "true";
defparam \rfile[31][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N8
cycloneive_lcell_comb \rfile[23][11]~feeder (
// Equation(s):
// \rfile[23][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[23][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[23][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[23][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N9
dffeas \rfile[23][11] (
	.clk(!CLK),
	.d(\rfile[23][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][11] .is_wysiwyg = "true";
defparam \rfile[23][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N6
cycloneive_lcell_comb \rfile[19][11]~feeder (
// Equation(s):
// \rfile[19][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[19][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[19][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[19][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N7
dffeas \rfile[19][11] (
	.clk(!CLK),
	.d(\rfile[19][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][11] .is_wysiwyg = "true";
defparam \rfile[19][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N20
cycloneive_lcell_comb \Mux52~7 (
// Equation(s):
// \Mux52~7_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[23][11]~q )) # (!instruction_D[18] & ((\rfile[19][11]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[23][11]~q ),
	.datad(\rfile[19][11]~q ),
	.cin(gnd),
	.combout(\Mux52~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~7 .lut_mask = 16'hD9C8;
defparam \Mux52~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y28_N26
cycloneive_lcell_comb \Mux52~8 (
// Equation(s):
// \Mux52~8_combout  = (instruction_D[19] & ((\Mux52~7_combout  & ((\rfile[31][11]~q ))) # (!\Mux52~7_combout  & (\rfile[27][11]~q )))) # (!instruction_D[19] & (((\Mux52~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[27][11]~q ),
	.datac(\rfile[31][11]~q ),
	.datad(\Mux52~7_combout ),
	.cin(gnd),
	.combout(\Mux52~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~8 .lut_mask = 16'hF588;
defparam \Mux52~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y29_N2
cycloneive_lcell_comb \rfile[29][11]~feeder (
// Equation(s):
// \rfile[29][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[29][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[29][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[29][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X77_Y29_N3
dffeas \rfile[29][11] (
	.clk(!CLK),
	.d(\rfile[29][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][11] .is_wysiwyg = "true";
defparam \rfile[29][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y30_N11
dffeas \rfile[17][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][11] .is_wysiwyg = "true";
defparam \rfile[17][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y30_N1
dffeas \rfile[21][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][11] .is_wysiwyg = "true";
defparam \rfile[21][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N10
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[21][11]~q )))) # (!instruction_D[18] & (!instruction_D[19] & (\rfile[17][11]~q )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[17][11]~q ),
	.datad(\rfile[21][11]~q ),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'hBA98;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y29_N12
cycloneive_lcell_comb \rfile[25][11]~feeder (
// Equation(s):
// \rfile[25][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[25][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[25][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[25][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X77_Y29_N13
dffeas \rfile[25][11] (
	.clk(!CLK),
	.d(\rfile[25][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][11] .is_wysiwyg = "true";
defparam \rfile[25][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X77_Y29_N24
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (instruction_D[19] & ((\Mux52~0_combout  & (\rfile[29][11]~q )) # (!\Mux52~0_combout  & ((\rfile[25][11]~q ))))) # (!instruction_D[19] & (((\Mux52~0_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[29][11]~q ),
	.datac(\Mux52~0_combout ),
	.datad(\rfile[25][11]~q ),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hDAD0;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N8
cycloneive_lcell_comb \rfile[18][11]~feeder (
// Equation(s):
// \rfile[18][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[18][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[18][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[18][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N9
dffeas \rfile[18][11] (
	.clk(!CLK),
	.d(\rfile[18][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][11] .is_wysiwyg = "true";
defparam \rfile[18][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N4
cycloneive_lcell_comb \Mux52~2 (
// Equation(s):
// \Mux52~2_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[26][11]~q )) # (!instruction_D[19] & ((\rfile[18][11]~q )))))

	.dataa(\rfile[26][11]~q ),
	.datab(instruction_D_18),
	.datac(instruction_D_19),
	.datad(\rfile[18][11]~q ),
	.cin(gnd),
	.combout(\Mux52~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~2 .lut_mask = 16'hE3E0;
defparam \Mux52~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N10
cycloneive_lcell_comb \rfile[22][11]~feeder (
// Equation(s):
// \rfile[22][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[22][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[22][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[22][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N11
dffeas \rfile[22][11] (
	.clk(!CLK),
	.d(\rfile[22][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][11] .is_wysiwyg = "true";
defparam \rfile[22][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N4
cycloneive_lcell_comb \Mux52~3 (
// Equation(s):
// \Mux52~3_combout  = (instruction_D[18] & ((\Mux52~2_combout  & (\rfile[30][11]~q )) # (!\Mux52~2_combout  & ((\rfile[22][11]~q ))))) # (!instruction_D[18] & (((\Mux52~2_combout ))))

	.dataa(\rfile[30][11]~q ),
	.datab(instruction_D_18),
	.datac(\Mux52~2_combout ),
	.datad(\rfile[22][11]~q ),
	.cin(gnd),
	.combout(\Mux52~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~3 .lut_mask = 16'hBCB0;
defparam \Mux52~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N18
cycloneive_lcell_comb \rfile[20][11]~feeder (
// Equation(s):
// \rfile[20][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[20][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[20][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[20][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N19
dffeas \rfile[20][11] (
	.clk(!CLK),
	.d(\rfile[20][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][11] .is_wysiwyg = "true";
defparam \rfile[20][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N15
dffeas \rfile[24][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][11] .is_wysiwyg = "true";
defparam \rfile[24][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N21
dffeas \rfile[16][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][11] .is_wysiwyg = "true";
defparam \rfile[16][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N20
cycloneive_lcell_comb \Mux52~4 (
// Equation(s):
// \Mux52~4_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[24][11]~q )) # (!instruction_D[19] & ((\rfile[16][11]~q )))))

	.dataa(instruction_D_18),
	.datab(\rfile[24][11]~q ),
	.datac(\rfile[16][11]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux52~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~4 .lut_mask = 16'hEE50;
defparam \Mux52~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y32_N25
dffeas \rfile[28][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][11] .is_wysiwyg = "true";
defparam \rfile[28][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N16
cycloneive_lcell_comb \Mux52~5 (
// Equation(s):
// \Mux52~5_combout  = (instruction_D[18] & ((\Mux52~4_combout  & ((\rfile[28][11]~q ))) # (!\Mux52~4_combout  & (\rfile[20][11]~q )))) # (!instruction_D[18] & (((\Mux52~4_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[20][11]~q ),
	.datac(\Mux52~4_combout ),
	.datad(\rfile[28][11]~q ),
	.cin(gnd),
	.combout(\Mux52~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~5 .lut_mask = 16'hF858;
defparam \Mux52~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N14
cycloneive_lcell_comb \Mux52~6 (
// Equation(s):
// \Mux52~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux52~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & ((\Mux52~5_combout ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux52~3_combout ),
	.datad(\Mux52~5_combout ),
	.cin(gnd),
	.combout(\Mux52~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~6 .lut_mask = 16'hB9A8;
defparam \Mux52~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N31
dffeas \rfile[15][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][11] .is_wysiwyg = "true";
defparam \rfile[15][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N12
cycloneive_lcell_comb \rfile[14][11]~feeder (
// Equation(s):
// \rfile[14][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[14][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[14][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N13
dffeas \rfile[14][11] (
	.clk(!CLK),
	.d(\rfile[14][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][11] .is_wysiwyg = "true";
defparam \rfile[14][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N11
dffeas \rfile[12][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][11] .is_wysiwyg = "true";
defparam \rfile[12][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N22
cycloneive_lcell_comb \rfile[13][11]~feeder (
// Equation(s):
// \rfile[13][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[13][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[13][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[13][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N23
dffeas \rfile[13][11] (
	.clk(!CLK),
	.d(\rfile[13][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][11] .is_wysiwyg = "true";
defparam \rfile[13][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N10
cycloneive_lcell_comb \Mux52~17 (
// Equation(s):
// \Mux52~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][11]~q ))) # (!instruction_D[16] & (\rfile[12][11]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][11]~q ),
	.datad(\rfile[13][11]~q ),
	.cin(gnd),
	.combout(\Mux52~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~17 .lut_mask = 16'hDC98;
defparam \Mux52~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N28
cycloneive_lcell_comb \Mux52~18 (
// Equation(s):
// \Mux52~18_combout  = (instruction_D[17] & ((\Mux52~17_combout  & (\rfile[15][11]~q )) # (!\Mux52~17_combout  & ((\rfile[14][11]~q ))))) # (!instruction_D[17] & (((\Mux52~17_combout ))))

	.dataa(\rfile[15][11]~q ),
	.datab(\rfile[14][11]~q ),
	.datac(instruction_D_17),
	.datad(\Mux52~17_combout ),
	.cin(gnd),
	.combout(\Mux52~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~18 .lut_mask = 16'hAFC0;
defparam \Mux52~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N21
dffeas \rfile[7][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][11] .is_wysiwyg = "true";
defparam \rfile[7][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N5
dffeas \rfile[4][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][11] .is_wysiwyg = "true";
defparam \rfile[4][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N15
dffeas \rfile[5][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][11] .is_wysiwyg = "true";
defparam \rfile[5][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N4
cycloneive_lcell_comb \Mux52~12 (
// Equation(s):
// \Mux52~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][11]~q ))) # (!instruction_D[16] & (\rfile[4][11]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][11]~q ),
	.datad(\rfile[5][11]~q ),
	.cin(gnd),
	.combout(\Mux52~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~12 .lut_mask = 16'hDC98;
defparam \Mux52~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N20
cycloneive_lcell_comb \Mux52~13 (
// Equation(s):
// \Mux52~13_combout  = (instruction_D[17] & ((\Mux52~12_combout  & ((\rfile[7][11]~q ))) # (!\Mux52~12_combout  & (\rfile[6][11]~q )))) # (!instruction_D[17] & (((\Mux52~12_combout ))))

	.dataa(\rfile[6][11]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[7][11]~q ),
	.datad(\Mux52~12_combout ),
	.cin(gnd),
	.combout(\Mux52~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~13 .lut_mask = 16'hF388;
defparam \Mux52~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N15
dffeas \rfile[2][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][11] .is_wysiwyg = "true";
defparam \rfile[2][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N15
dffeas \rfile[1][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][11] .is_wysiwyg = "true";
defparam \rfile[1][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N12
cycloneive_lcell_comb \rfile[3][11]~feeder (
// Equation(s):
// \rfile[3][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_11),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[3][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[3][11]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[3][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y27_N13
dffeas \rfile[3][11] (
	.clk(!CLK),
	.d(\rfile[3][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][11] .is_wysiwyg = "true";
defparam \rfile[3][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N14
cycloneive_lcell_comb \Mux52~14 (
// Equation(s):
// \Mux52~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][11]~q ))) # (!instruction_D[17] & (\rfile[1][11]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[1][11]~q ),
	.datad(\rfile[3][11]~q ),
	.cin(gnd),
	.combout(\Mux52~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~14 .lut_mask = 16'hA820;
defparam \Mux52~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N24
cycloneive_lcell_comb \Mux52~15 (
// Equation(s):
// \Mux52~15_combout  = (\Mux52~14_combout ) # ((instruction_D[17] & (!instruction_D[16] & \rfile[2][11]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[2][11]~q ),
	.datad(\Mux52~14_combout ),
	.cin(gnd),
	.combout(\Mux52~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~15 .lut_mask = 16'hFF20;
defparam \Mux52~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N22
cycloneive_lcell_comb \Mux52~16 (
// Equation(s):
// \Mux52~16_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\Mux52~13_combout )) # (!instruction_D[18] & ((\Mux52~15_combout )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux52~13_combout ),
	.datad(\Mux52~15_combout ),
	.cin(gnd),
	.combout(\Mux52~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~16 .lut_mask = 16'hD9C8;
defparam \Mux52~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N14
cycloneive_lcell_comb \rfile[9][11]~feeder (
// Equation(s):
// \rfile[9][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_11),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[9][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][11]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[9][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N15
dffeas \rfile[9][11] (
	.clk(!CLK),
	.d(\rfile[9][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][11] .is_wysiwyg = "true";
defparam \rfile[9][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y35_N25
dffeas \rfile[11][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][11] .is_wysiwyg = "true";
defparam \rfile[11][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N25
dffeas \rfile[10][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][11] .is_wysiwyg = "true";
defparam \rfile[10][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N7
dffeas \rfile[8][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][11] .is_wysiwyg = "true";
defparam \rfile[8][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N24
cycloneive_lcell_comb \Mux52~10 (
// Equation(s):
// \Mux52~10_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\rfile[10][11]~q )) # (!instruction_D[17] & ((\rfile[8][11]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[10][11]~q ),
	.datad(\rfile[8][11]~q ),
	.cin(gnd),
	.combout(\Mux52~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~10 .lut_mask = 16'hD9C8;
defparam \Mux52~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N24
cycloneive_lcell_comb \Mux52~11 (
// Equation(s):
// \Mux52~11_combout  = (instruction_D[16] & ((\Mux52~10_combout  & ((\rfile[11][11]~q ))) # (!\Mux52~10_combout  & (\rfile[9][11]~q )))) # (!instruction_D[16] & (((\Mux52~10_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[9][11]~q ),
	.datac(\rfile[11][11]~q ),
	.datad(\Mux52~10_combout ),
	.cin(gnd),
	.combout(\Mux52~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~11 .lut_mask = 16'hF588;
defparam \Mux52~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N23
dffeas \rfile[25][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][10] .is_wysiwyg = "true";
defparam \rfile[25][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N22
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (instruction_D[19] & (((\rfile[25][10]~q ) # (instruction_D[18])))) # (!instruction_D[19] & (\rfile[17][10]~q  & ((!instruction_D[18]))))

	.dataa(\rfile[17][10]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[25][10]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'hCCE2;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N9
dffeas \rfile[21][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][10] .is_wysiwyg = "true";
defparam \rfile[21][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y28_N12
cycloneive_lcell_comb \rfile[29][10]~feeder (
// Equation(s):
// \rfile[29][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_10),
	.cin(gnd),
	.combout(\rfile[29][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[29][10]~feeder .lut_mask = 16'hFF00;
defparam \rfile[29][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y28_N13
dffeas \rfile[29][10] (
	.clk(!CLK),
	.d(\rfile[29][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][10] .is_wysiwyg = "true";
defparam \rfile[29][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N12
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (instruction_D[18] & ((\Mux53~0_combout  & ((\rfile[29][10]~q ))) # (!\Mux53~0_combout  & (\rfile[21][10]~q )))) # (!instruction_D[18] & (\Mux53~0_combout ))

	.dataa(instruction_D_18),
	.datab(\Mux53~0_combout ),
	.datac(\rfile[21][10]~q ),
	.datad(\rfile[29][10]~q ),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'hEC64;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N26
cycloneive_lcell_comb \rfile[23][10]~feeder (
// Equation(s):
// \rfile[23][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_10),
	.cin(gnd),
	.combout(\rfile[23][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[23][10]~feeder .lut_mask = 16'hFF00;
defparam \rfile[23][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N27
dffeas \rfile[23][10] (
	.clk(!CLK),
	.d(\rfile[23][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][10] .is_wysiwyg = "true";
defparam \rfile[23][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y28_N23
dffeas \rfile[31][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][10] .is_wysiwyg = "true";
defparam \rfile[31][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y28_N22
cycloneive_lcell_comb \rfile[27][10]~feeder (
// Equation(s):
// \rfile[27][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_10),
	.cin(gnd),
	.combout(\rfile[27][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[27][10]~feeder .lut_mask = 16'hFF00;
defparam \rfile[27][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y28_N23
dffeas \rfile[27][10] (
	.clk(!CLK),
	.d(\rfile[27][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][10] .is_wysiwyg = "true";
defparam \rfile[27][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N8
cycloneive_lcell_comb \rfile[19][10]~feeder (
// Equation(s):
// \rfile[19][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_10),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[19][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[19][10]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[19][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y28_N9
dffeas \rfile[19][10] (
	.clk(!CLK),
	.d(\rfile[19][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][10] .is_wysiwyg = "true";
defparam \rfile[19][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y28_N20
cycloneive_lcell_comb \Mux53~7 (
// Equation(s):
// \Mux53~7_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[27][10]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[19][10]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[27][10]~q ),
	.datad(\rfile[19][10]~q ),
	.cin(gnd),
	.combout(\Mux53~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~7 .lut_mask = 16'hB9A8;
defparam \Mux53~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N24
cycloneive_lcell_comb \Mux53~8 (
// Equation(s):
// \Mux53~8_combout  = (instruction_D[18] & ((\Mux53~7_combout  & ((\rfile[31][10]~q ))) # (!\Mux53~7_combout  & (\rfile[23][10]~q )))) # (!instruction_D[18] & (((\Mux53~7_combout ))))

	.dataa(\rfile[23][10]~q ),
	.datab(\rfile[31][10]~q ),
	.datac(instruction_D_18),
	.datad(\Mux53~7_combout ),
	.cin(gnd),
	.combout(\Mux53~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~8 .lut_mask = 16'hCFA0;
defparam \Mux53~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y32_N5
dffeas \rfile[28][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][10] .is_wysiwyg = "true";
defparam \rfile[28][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N6
cycloneive_lcell_comb \rfile[24][10]~feeder (
// Equation(s):
// \rfile[24][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_10),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[24][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[24][10]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[24][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y32_N7
dffeas \rfile[24][10] (
	.clk(!CLK),
	.d(\rfile[24][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][10] .is_wysiwyg = "true";
defparam \rfile[24][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N21
dffeas \rfile[20][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][10] .is_wysiwyg = "true";
defparam \rfile[20][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N27
dffeas \rfile[16][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][10] .is_wysiwyg = "true";
defparam \rfile[16][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N20
cycloneive_lcell_comb \Mux53~4 (
// Equation(s):
// \Mux53~4_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[20][10]~q )) # (!instruction_D[18] & ((\rfile[16][10]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[20][10]~q ),
	.datad(\rfile[16][10]~q ),
	.cin(gnd),
	.combout(\Mux53~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~4 .lut_mask = 16'hD9C8;
defparam \Mux53~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N30
cycloneive_lcell_comb \Mux53~5 (
// Equation(s):
// \Mux53~5_combout  = (instruction_D[19] & ((\Mux53~4_combout  & (\rfile[28][10]~q )) # (!\Mux53~4_combout  & ((\rfile[24][10]~q ))))) # (!instruction_D[19] & (((\Mux53~4_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[28][10]~q ),
	.datac(\rfile[24][10]~q ),
	.datad(\Mux53~4_combout ),
	.cin(gnd),
	.combout(\Mux53~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~5 .lut_mask = 16'hDDA0;
defparam \Mux53~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y36_N21
dffeas \rfile[30][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][10] .is_wysiwyg = "true";
defparam \rfile[30][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y36_N26
cycloneive_lcell_comb \rfile[18][10]~feeder (
// Equation(s):
// \rfile[18][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_10),
	.cin(gnd),
	.combout(\rfile[18][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[18][10]~feeder .lut_mask = 16'hFF00;
defparam \rfile[18][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y36_N27
dffeas \rfile[18][10] (
	.clk(!CLK),
	.d(\rfile[18][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][10] .is_wysiwyg = "true";
defparam \rfile[18][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y36_N12
cycloneive_lcell_comb \rfile[22][10]~feeder (
// Equation(s):
// \rfile[22][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_10),
	.cin(gnd),
	.combout(\rfile[22][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[22][10]~feeder .lut_mask = 16'hFF00;
defparam \rfile[22][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y36_N13
dffeas \rfile[22][10] (
	.clk(!CLK),
	.d(\rfile[22][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][10] .is_wysiwyg = "true";
defparam \rfile[22][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y36_N24
cycloneive_lcell_comb \Mux53~2 (
// Equation(s):
// \Mux53~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[22][10]~q ))) # (!instruction_D[18] & (\rfile[18][10]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][10]~q ),
	.datad(\rfile[22][10]~q ),
	.cin(gnd),
	.combout(\Mux53~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~2 .lut_mask = 16'hDC98;
defparam \Mux53~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N20
cycloneive_lcell_comb \Mux53~3 (
// Equation(s):
// \Mux53~3_combout  = (instruction_D[19] & ((\Mux53~2_combout  & ((\rfile[30][10]~q ))) # (!\Mux53~2_combout  & (\rfile[26][10]~q )))) # (!instruction_D[19] & (((\Mux53~2_combout ))))

	.dataa(\rfile[26][10]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[30][10]~q ),
	.datad(\Mux53~2_combout ),
	.cin(gnd),
	.combout(\Mux53~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~3 .lut_mask = 16'hF388;
defparam \Mux53~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N28
cycloneive_lcell_comb \Mux53~6 (
// Equation(s):
// \Mux53~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux53~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & (\Mux53~5_combout )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux53~5_combout ),
	.datad(\Mux53~3_combout ),
	.cin(gnd),
	.combout(\Mux53~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~6 .lut_mask = 16'hBA98;
defparam \Mux53~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N21
dffeas \rfile[6][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][10] .is_wysiwyg = "true";
defparam \rfile[6][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y28_N19
dffeas \rfile[7][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][10] .is_wysiwyg = "true";
defparam \rfile[7][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y28_N21
dffeas \rfile[4][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][10] .is_wysiwyg = "true";
defparam \rfile[4][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N9
dffeas \rfile[5][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][10] .is_wysiwyg = "true";
defparam \rfile[5][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N20
cycloneive_lcell_comb \Mux53~10 (
// Equation(s):
// \Mux53~10_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][10]~q ))) # (!instruction_D[16] & (\rfile[4][10]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][10]~q ),
	.datad(\rfile[5][10]~q ),
	.cin(gnd),
	.combout(\Mux53~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~10 .lut_mask = 16'hDC98;
defparam \Mux53~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N18
cycloneive_lcell_comb \Mux53~11 (
// Equation(s):
// \Mux53~11_combout  = (instruction_D[17] & ((\Mux53~10_combout  & ((\rfile[7][10]~q ))) # (!\Mux53~10_combout  & (\rfile[6][10]~q )))) # (!instruction_D[17] & (((\Mux53~10_combout ))))

	.dataa(\rfile[6][10]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[7][10]~q ),
	.datad(\Mux53~10_combout ),
	.cin(gnd),
	.combout(\Mux53~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~11 .lut_mask = 16'hF388;
defparam \Mux53~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N11
dffeas \rfile[15][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][10] .is_wysiwyg = "true";
defparam \rfile[15][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N2
cycloneive_lcell_comb \rfile[14][10]~feeder (
// Equation(s):
// \rfile[14][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_10),
	.cin(gnd),
	.combout(\rfile[14][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][10]~feeder .lut_mask = 16'hFF00;
defparam \rfile[14][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N3
dffeas \rfile[14][10] (
	.clk(!CLK),
	.d(\rfile[14][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][10] .is_wysiwyg = "true";
defparam \rfile[14][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N8
cycloneive_lcell_comb \rfile[13][10]~feeder (
// Equation(s):
// \rfile[13][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_10),
	.cin(gnd),
	.combout(\rfile[13][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[13][10]~feeder .lut_mask = 16'hFF00;
defparam \rfile[13][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N9
dffeas \rfile[13][10] (
	.clk(!CLK),
	.d(\rfile[13][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][10] .is_wysiwyg = "true";
defparam \rfile[13][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N19
dffeas \rfile[12][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][10] .is_wysiwyg = "true";
defparam \rfile[12][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N30
cycloneive_lcell_comb \Mux53~17 (
// Equation(s):
// \Mux53~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][10]~q )))) # (!instruction_D[16] & (!instruction_D[17] & ((\rfile[12][10]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[13][10]~q ),
	.datad(\rfile[12][10]~q ),
	.cin(gnd),
	.combout(\Mux53~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~17 .lut_mask = 16'hB9A8;
defparam \Mux53~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N14
cycloneive_lcell_comb \Mux53~18 (
// Equation(s):
// \Mux53~18_combout  = (instruction_D[17] & ((\Mux53~17_combout  & (\rfile[15][10]~q )) # (!\Mux53~17_combout  & ((\rfile[14][10]~q ))))) # (!instruction_D[17] & (((\Mux53~17_combout ))))

	.dataa(\rfile[15][10]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[14][10]~q ),
	.datad(\Mux53~17_combout ),
	.cin(gnd),
	.combout(\Mux53~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~18 .lut_mask = 16'hBBC0;
defparam \Mux53~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N28
cycloneive_lcell_comb \rfile[11][10]~feeder (
// Equation(s):
// \rfile[11][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_10),
	.cin(gnd),
	.combout(\rfile[11][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][10]~feeder .lut_mask = 16'hFF00;
defparam \rfile[11][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y27_N29
dffeas \rfile[11][10] (
	.clk(!CLK),
	.d(\rfile[11][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][10] .is_wysiwyg = "true";
defparam \rfile[11][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N12
cycloneive_lcell_comb \rfile[9][10]~feeder (
// Equation(s):
// \rfile[9][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_10),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[9][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][10]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[9][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N13
dffeas \rfile[9][10] (
	.clk(!CLK),
	.d(\rfile[9][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][10] .is_wysiwyg = "true";
defparam \rfile[9][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N27
dffeas \rfile[8][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][10] .is_wysiwyg = "true";
defparam \rfile[8][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N29
dffeas \rfile[10][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][10] .is_wysiwyg = "true";
defparam \rfile[10][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N26
cycloneive_lcell_comb \Mux53~12 (
// Equation(s):
// \Mux53~12_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][10]~q ))) # (!instruction_D[17] & (\rfile[8][10]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[8][10]~q ),
	.datad(\rfile[10][10]~q ),
	.cin(gnd),
	.combout(\Mux53~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~12 .lut_mask = 16'hDC98;
defparam \Mux53~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N18
cycloneive_lcell_comb \Mux53~13 (
// Equation(s):
// \Mux53~13_combout  = (instruction_D[16] & ((\Mux53~12_combout  & (\rfile[11][10]~q )) # (!\Mux53~12_combout  & ((\rfile[9][10]~q ))))) # (!instruction_D[16] & (((\Mux53~12_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][10]~q ),
	.datac(\rfile[9][10]~q ),
	.datad(\Mux53~12_combout ),
	.cin(gnd),
	.combout(\Mux53~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~13 .lut_mask = 16'hDDA0;
defparam \Mux53~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N4
cycloneive_lcell_comb \rfile[2][10]~feeder (
// Equation(s):
// \rfile[2][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_10),
	.cin(gnd),
	.combout(\rfile[2][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][10]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y27_N5
dffeas \rfile[2][10] (
	.clk(!CLK),
	.d(\rfile[2][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][10] .is_wysiwyg = "true";
defparam \rfile[2][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N30
cycloneive_lcell_comb \rfile[3][10]~feeder (
// Equation(s):
// \rfile[3][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_10),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[3][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[3][10]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[3][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N31
dffeas \rfile[3][10] (
	.clk(!CLK),
	.d(\rfile[3][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][10] .is_wysiwyg = "true";
defparam \rfile[3][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N24
cycloneive_lcell_comb \rfile[1][10]~feeder (
// Equation(s):
// \rfile[1][10]~feeder_combout  = \wdat_WB[10]~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_10),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[1][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[1][10]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[1][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N25
dffeas \rfile[1][10] (
	.clk(!CLK),
	.d(\rfile[1][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][10] .is_wysiwyg = "true";
defparam \rfile[1][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N6
cycloneive_lcell_comb \Mux53~14 (
// Equation(s):
// \Mux53~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][10]~q )) # (!instruction_D[17] & ((\rfile[1][10]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[3][10]~q ),
	.datad(\rfile[1][10]~q ),
	.cin(gnd),
	.combout(\Mux53~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~14 .lut_mask = 16'hA280;
defparam \Mux53~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N2
cycloneive_lcell_comb \Mux53~15 (
// Equation(s):
// \Mux53~15_combout  = (\Mux53~14_combout ) # ((!instruction_D[16] & (instruction_D[17] & \rfile[2][10]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[2][10]~q ),
	.datad(\Mux53~14_combout ),
	.cin(gnd),
	.combout(\Mux53~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~15 .lut_mask = 16'hFF40;
defparam \Mux53~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N0
cycloneive_lcell_comb \Mux53~16 (
// Equation(s):
// \Mux53~16_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & (\Mux53~13_combout )) # (!instruction_D[19] & ((\Mux53~15_combout )))))

	.dataa(instruction_D_18),
	.datab(\Mux53~13_combout ),
	.datac(instruction_D_19),
	.datad(\Mux53~15_combout ),
	.cin(gnd),
	.combout(\Mux53~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~16 .lut_mask = 16'hE5E0;
defparam \Mux53~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N30
cycloneive_lcell_comb \rfile[17][7]~feeder (
// Equation(s):
// \rfile[17][7]~feeder_combout  = \wdat_WB[7]~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[17][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[17][7]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[17][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y28_N31
dffeas \rfile[17][7] (
	.clk(!CLK),
	.d(\rfile[17][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][7] .is_wysiwyg = "true";
defparam \rfile[17][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N9
dffeas \rfile[21][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][7] .is_wysiwyg = "true";
defparam \rfile[21][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N18
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[21][7]~q ))) # (!instruction_D[18] & (\rfile[17][7]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[17][7]~q ),
	.datad(\rfile[21][7]~q ),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'hDC98;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N1
dffeas \rfile[29][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][7] .is_wysiwyg = "true";
defparam \rfile[29][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N17
dffeas \rfile[25][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][7] .is_wysiwyg = "true";
defparam \rfile[25][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N0
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (instruction_D[19] & ((\Mux56~0_combout  & (\rfile[29][7]~q )) # (!\Mux56~0_combout  & ((\rfile[25][7]~q ))))) # (!instruction_D[19] & (\Mux56~0_combout ))

	.dataa(instruction_D_19),
	.datab(\Mux56~0_combout ),
	.datac(\rfile[29][7]~q ),
	.datad(\rfile[25][7]~q ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hE6C4;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y29_N25
dffeas \rfile[31][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][7] .is_wysiwyg = "true";
defparam \rfile[31][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N31
dffeas \rfile[27][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][7] .is_wysiwyg = "true";
defparam \rfile[27][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N15
dffeas \rfile[19][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][7] .is_wysiwyg = "true";
defparam \rfile[19][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N17
dffeas \rfile[23][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][7] .is_wysiwyg = "true";
defparam \rfile[23][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N14
cycloneive_lcell_comb \Mux56~7 (
// Equation(s):
// \Mux56~7_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[23][7]~q ))) # (!instruction_D[18] & (\rfile[19][7]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[19][7]~q ),
	.datad(\rfile[23][7]~q ),
	.cin(gnd),
	.combout(\Mux56~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~7 .lut_mask = 16'hDC98;
defparam \Mux56~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N30
cycloneive_lcell_comb \Mux56~8 (
// Equation(s):
// \Mux56~8_combout  = (instruction_D[19] & ((\Mux56~7_combout  & (\rfile[31][7]~q )) # (!\Mux56~7_combout  & ((\rfile[27][7]~q ))))) # (!instruction_D[19] & (((\Mux56~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[31][7]~q ),
	.datac(\rfile[27][7]~q ),
	.datad(\Mux56~7_combout ),
	.cin(gnd),
	.combout(\Mux56~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~8 .lut_mask = 16'hDDA0;
defparam \Mux56~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N22
cycloneive_lcell_comb \rfile[28][7]~feeder (
// Equation(s):
// \rfile[28][7]~feeder_combout  = \wdat_WB[7]~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_7),
	.cin(gnd),
	.combout(\rfile[28][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][7]~feeder .lut_mask = 16'hFF00;
defparam \rfile[28][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y32_N23
dffeas \rfile[28][7] (
	.clk(!CLK),
	.d(\rfile[28][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][7] .is_wysiwyg = "true";
defparam \rfile[28][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y32_N23
dffeas \rfile[20][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][7] .is_wysiwyg = "true";
defparam \rfile[20][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N30
cycloneive_lcell_comb \rfile[24][7]~feeder (
// Equation(s):
// \rfile[24][7]~feeder_combout  = \wdat_WB[7]~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_7),
	.cin(gnd),
	.combout(\rfile[24][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[24][7]~feeder .lut_mask = 16'hFF00;
defparam \rfile[24][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y32_N31
dffeas \rfile[24][7] (
	.clk(!CLK),
	.d(\rfile[24][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][7] .is_wysiwyg = "true";
defparam \rfile[24][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N16
cycloneive_lcell_comb \rfile[16][7]~feeder (
// Equation(s):
// \rfile[16][7]~feeder_combout  = \wdat_WB[7]~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[16][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[16][7]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[16][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y32_N17
dffeas \rfile[16][7] (
	.clk(!CLK),
	.d(\rfile[16][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][7] .is_wysiwyg = "true";
defparam \rfile[16][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N8
cycloneive_lcell_comb \Mux56~4 (
// Equation(s):
// \Mux56~4_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[24][7]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[16][7]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[24][7]~q ),
	.datad(\rfile[16][7]~q ),
	.cin(gnd),
	.combout(\Mux56~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~4 .lut_mask = 16'hB9A8;
defparam \Mux56~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N22
cycloneive_lcell_comb \Mux56~5 (
// Equation(s):
// \Mux56~5_combout  = (instruction_D[18] & ((\Mux56~4_combout  & (\rfile[28][7]~q )) # (!\Mux56~4_combout  & ((\rfile[20][7]~q ))))) # (!instruction_D[18] & (((\Mux56~4_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[28][7]~q ),
	.datac(\rfile[20][7]~q ),
	.datad(\Mux56~4_combout ),
	.cin(gnd),
	.combout(\Mux56~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~5 .lut_mask = 16'hDDA0;
defparam \Mux56~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y35_N21
dffeas \rfile[22][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][7] .is_wysiwyg = "true";
defparam \rfile[22][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y35_N7
dffeas \rfile[30][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][7] .is_wysiwyg = "true";
defparam \rfile[30][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N30
cycloneive_lcell_comb \rfile[26][7]~feeder (
// Equation(s):
// \rfile[26][7]~feeder_combout  = \wdat_WB[7]~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_7),
	.cin(gnd),
	.combout(\rfile[26][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[26][7]~feeder .lut_mask = 16'hFF00;
defparam \rfile[26][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y36_N31
dffeas \rfile[26][7] (
	.clk(!CLK),
	.d(\rfile[26][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][7] .is_wysiwyg = "true";
defparam \rfile[26][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N6
cycloneive_lcell_comb \rfile[18][7]~feeder (
// Equation(s):
// \rfile[18][7]~feeder_combout  = \wdat_WB[7]~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[18][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[18][7]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[18][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y35_N7
dffeas \rfile[18][7] (
	.clk(!CLK),
	.d(\rfile[18][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][7] .is_wysiwyg = "true";
defparam \rfile[18][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N4
cycloneive_lcell_comb \Mux56~2 (
// Equation(s):
// \Mux56~2_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[26][7]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[18][7]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[26][7]~q ),
	.datad(\rfile[18][7]~q ),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~2 .lut_mask = 16'hB9A8;
defparam \Mux56~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N6
cycloneive_lcell_comb \Mux56~3 (
// Equation(s):
// \Mux56~3_combout  = (instruction_D[18] & ((\Mux56~2_combout  & ((\rfile[30][7]~q ))) # (!\Mux56~2_combout  & (\rfile[22][7]~q )))) # (!instruction_D[18] & (((\Mux56~2_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[22][7]~q ),
	.datac(\rfile[30][7]~q ),
	.datad(\Mux56~2_combout ),
	.cin(gnd),
	.combout(\Mux56~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~3 .lut_mask = 16'hF588;
defparam \Mux56~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N6
cycloneive_lcell_comb \Mux56~6 (
// Equation(s):
// \Mux56~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux56~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & (\Mux56~5_combout )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux56~5_combout ),
	.datad(\Mux56~3_combout ),
	.cin(gnd),
	.combout(\Mux56~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~6 .lut_mask = 16'hBA98;
defparam \Mux56~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N8
cycloneive_lcell_comb \rfile[15][7]~feeder (
// Equation(s):
// \rfile[15][7]~feeder_combout  = \wdat_WB[7]~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_7),
	.cin(gnd),
	.combout(\rfile[15][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][7]~feeder .lut_mask = 16'hFF00;
defparam \rfile[15][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N9
dffeas \rfile[15][7] (
	.clk(!CLK),
	.d(\rfile[15][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][7] .is_wysiwyg = "true";
defparam \rfile[15][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y33_N5
dffeas \rfile[14][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][7] .is_wysiwyg = "true";
defparam \rfile[14][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N17
dffeas \rfile[13][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][7] .is_wysiwyg = "true";
defparam \rfile[13][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N16
cycloneive_lcell_comb \Mux56~17 (
// Equation(s):
// \Mux56~17_combout  = (instruction_D[16] & (((\rfile[13][7]~q ) # (instruction_D[17])))) # (!instruction_D[16] & (\rfile[12][7]~q  & ((!instruction_D[17]))))

	.dataa(\rfile[12][7]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[13][7]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux56~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~17 .lut_mask = 16'hCCE2;
defparam \Mux56~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N2
cycloneive_lcell_comb \Mux56~18 (
// Equation(s):
// \Mux56~18_combout  = (instruction_D[17] & ((\Mux56~17_combout  & (\rfile[15][7]~q )) # (!\Mux56~17_combout  & ((\rfile[14][7]~q ))))) # (!instruction_D[17] & (((\Mux56~17_combout ))))

	.dataa(\rfile[15][7]~q ),
	.datab(\rfile[14][7]~q ),
	.datac(instruction_D_17),
	.datad(\Mux56~17_combout ),
	.cin(gnd),
	.combout(\Mux56~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~18 .lut_mask = 16'hAFC0;
defparam \Mux56~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y28_N15
dffeas \rfile[4][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][7] .is_wysiwyg = "true";
defparam \rfile[4][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N21
dffeas \rfile[5][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][7] .is_wysiwyg = "true";
defparam \rfile[5][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N14
cycloneive_lcell_comb \Mux56~12 (
// Equation(s):
// \Mux56~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][7]~q ))) # (!instruction_D[16] & (\rfile[4][7]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][7]~q ),
	.datad(\rfile[5][7]~q ),
	.cin(gnd),
	.combout(\Mux56~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~12 .lut_mask = 16'hDC98;
defparam \Mux56~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N17
dffeas \rfile[7][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][7] .is_wysiwyg = "true";
defparam \rfile[7][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N8
cycloneive_lcell_comb \Mux56~13 (
// Equation(s):
// \Mux56~13_combout  = (\Mux56~12_combout  & (((\rfile[7][7]~q ) # (!instruction_D[17])))) # (!\Mux56~12_combout  & (\rfile[6][7]~q  & (instruction_D[17])))

	.dataa(\rfile[6][7]~q ),
	.datab(\Mux56~12_combout ),
	.datac(instruction_D_17),
	.datad(\rfile[7][7]~q ),
	.cin(gnd),
	.combout(\Mux56~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~13 .lut_mask = 16'hEC2C;
defparam \Mux56~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y27_N17
dffeas \rfile[3][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][7] .is_wysiwyg = "true";
defparam \rfile[3][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N7
dffeas \rfile[1][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][7] .is_wysiwyg = "true";
defparam \rfile[1][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N16
cycloneive_lcell_comb \Mux56~14 (
// Equation(s):
// \Mux56~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][7]~q )) # (!instruction_D[17] & ((\rfile[1][7]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[3][7]~q ),
	.datad(\rfile[1][7]~q ),
	.cin(gnd),
	.combout(\Mux56~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~14 .lut_mask = 16'hA280;
defparam \Mux56~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N0
cycloneive_lcell_comb \Mux56~15 (
// Equation(s):
// \Mux56~15_combout  = (\Mux56~14_combout ) # ((\rfile[2][7]~q  & (!instruction_D[16] & instruction_D[17])))

	.dataa(\rfile[2][7]~q ),
	.datab(instruction_D_16),
	.datac(instruction_D_17),
	.datad(\Mux56~14_combout ),
	.cin(gnd),
	.combout(\Mux56~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~15 .lut_mask = 16'hFF20;
defparam \Mux56~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N26
cycloneive_lcell_comb \Mux56~16 (
// Equation(s):
// \Mux56~16_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\Mux56~13_combout )) # (!instruction_D[18] & ((\Mux56~15_combout )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux56~13_combout ),
	.datad(\Mux56~15_combout ),
	.cin(gnd),
	.combout(\Mux56~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~16 .lut_mask = 16'hD9C8;
defparam \Mux56~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y35_N5
dffeas \rfile[10][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][7] .is_wysiwyg = "true";
defparam \rfile[10][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N19
dffeas \rfile[8][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][7] .is_wysiwyg = "true";
defparam \rfile[8][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N4
cycloneive_lcell_comb \Mux56~10 (
// Equation(s):
// \Mux56~10_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][7]~q )))) # (!instruction_D[17] & (!instruction_D[16] & ((\rfile[8][7]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[10][7]~q ),
	.datad(\rfile[8][7]~q ),
	.cin(gnd),
	.combout(\Mux56~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~10 .lut_mask = 16'hB9A8;
defparam \Mux56~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N1
dffeas \rfile[11][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][7] .is_wysiwyg = "true";
defparam \rfile[11][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N10
cycloneive_lcell_comb \rfile[9][7]~feeder (
// Equation(s):
// \rfile[9][7]~feeder_combout  = \wdat_WB[7]~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[9][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][7]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[9][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N11
dffeas \rfile[9][7] (
	.clk(!CLK),
	.d(\rfile[9][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][7] .is_wysiwyg = "true";
defparam \rfile[9][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N0
cycloneive_lcell_comb \Mux56~11 (
// Equation(s):
// \Mux56~11_combout  = (instruction_D[16] & ((\Mux56~10_combout  & (\rfile[11][7]~q )) # (!\Mux56~10_combout  & ((\rfile[9][7]~q ))))) # (!instruction_D[16] & (\Mux56~10_combout ))

	.dataa(instruction_D_16),
	.datab(\Mux56~10_combout ),
	.datac(\rfile[11][7]~q ),
	.datad(\rfile[9][7]~q ),
	.cin(gnd),
	.combout(\Mux56~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~11 .lut_mask = 16'hE6C4;
defparam \Mux56~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N2
cycloneive_lcell_comb \rfile[21][6]~feeder (
// Equation(s):
// \rfile[21][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[21][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][6]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[21][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N3
dffeas \rfile[21][6] (
	.clk(!CLK),
	.d(\rfile[21][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][6] .is_wysiwyg = "true";
defparam \rfile[21][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N6
cycloneive_lcell_comb \rfile[29][6]~feeder (
// Equation(s):
// \rfile[29][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_6),
	.cin(gnd),
	.combout(\rfile[29][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[29][6]~feeder .lut_mask = 16'hFF00;
defparam \rfile[29][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N7
dffeas \rfile[29][6] (
	.clk(!CLK),
	.d(\rfile[29][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][6] .is_wysiwyg = "true";
defparam \rfile[29][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N5
dffeas \rfile[25][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][6] .is_wysiwyg = "true";
defparam \rfile[25][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N7
dffeas \rfile[17][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][6] .is_wysiwyg = "true";
defparam \rfile[17][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N6
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (instruction_D[19] & ((\rfile[25][6]~q ) # ((instruction_D[18])))) # (!instruction_D[19] & (((\rfile[17][6]~q  & !instruction_D[18]))))

	.dataa(instruction_D_19),
	.datab(\rfile[25][6]~q ),
	.datac(\rfile[17][6]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'hAAD8;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N4
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (instruction_D[18] & ((\Mux57~0_combout  & ((\rfile[29][6]~q ))) # (!\Mux57~0_combout  & (\rfile[21][6]~q )))) # (!instruction_D[18] & (((\Mux57~0_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[21][6]~q ),
	.datac(\rfile[29][6]~q ),
	.datad(\Mux57~0_combout ),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hF588;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N21
dffeas \rfile[24][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][6] .is_wysiwyg = "true";
defparam \rfile[24][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y32_N19
dffeas \rfile[20][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][6] .is_wysiwyg = "true";
defparam \rfile[20][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y32_N29
dffeas \rfile[16][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][6] .is_wysiwyg = "true";
defparam \rfile[16][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N18
cycloneive_lcell_comb \Mux57~4 (
// Equation(s):
// \Mux57~4_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[20][6]~q )) # (!instruction_D[18] & ((\rfile[16][6]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[20][6]~q ),
	.datad(\rfile[16][6]~q ),
	.cin(gnd),
	.combout(\Mux57~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~4 .lut_mask = 16'hD9C8;
defparam \Mux57~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N18
cycloneive_lcell_comb \rfile[28][6]~feeder (
// Equation(s):
// \rfile[28][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[28][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][6]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[28][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N19
dffeas \rfile[28][6] (
	.clk(!CLK),
	.d(\rfile[28][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][6] .is_wysiwyg = "true";
defparam \rfile[28][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N30
cycloneive_lcell_comb \Mux57~5 (
// Equation(s):
// \Mux57~5_combout  = (instruction_D[19] & ((\Mux57~4_combout  & ((\rfile[28][6]~q ))) # (!\Mux57~4_combout  & (\rfile[24][6]~q )))) # (!instruction_D[19] & (((\Mux57~4_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[24][6]~q ),
	.datac(\Mux57~4_combout ),
	.datad(\rfile[28][6]~q ),
	.cin(gnd),
	.combout(\Mux57~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~5 .lut_mask = 16'hF858;
defparam \Mux57~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y35_N29
dffeas \rfile[30][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][6] .is_wysiwyg = "true";
defparam \rfile[30][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N4
cycloneive_lcell_comb \rfile[22][6]~feeder (
// Equation(s):
// \rfile[22][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[22][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[22][6]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[22][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y35_N5
dffeas \rfile[22][6] (
	.clk(!CLK),
	.d(\rfile[22][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][6] .is_wysiwyg = "true";
defparam \rfile[22][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N27
dffeas \rfile[18][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][6] .is_wysiwyg = "true";
defparam \rfile[18][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N10
cycloneive_lcell_comb \Mux57~2 (
// Equation(s):
// \Mux57~2_combout  = (instruction_D[19] & (((instruction_D[18])))) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[22][6]~q )) # (!instruction_D[18] & ((\rfile[18][6]~q )))))

	.dataa(instruction_D_19),
	.datab(\rfile[22][6]~q ),
	.datac(\rfile[18][6]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux57~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~2 .lut_mask = 16'hEE50;
defparam \Mux57~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N28
cycloneive_lcell_comb \Mux57~3 (
// Equation(s):
// \Mux57~3_combout  = (instruction_D[19] & ((\Mux57~2_combout  & ((\rfile[30][6]~q ))) # (!\Mux57~2_combout  & (\rfile[26][6]~q )))) # (!instruction_D[19] & (((\Mux57~2_combout ))))

	.dataa(\rfile[26][6]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[30][6]~q ),
	.datad(\Mux57~2_combout ),
	.cin(gnd),
	.combout(\Mux57~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~3 .lut_mask = 16'hF388;
defparam \Mux57~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N8
cycloneive_lcell_comb \Mux57~6 (
// Equation(s):
// \Mux57~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\Mux57~3_combout ))) # (!instruction_D[17] & (\Mux57~5_combout ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux57~5_combout ),
	.datad(\Mux57~3_combout ),
	.cin(gnd),
	.combout(\Mux57~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~6 .lut_mask = 16'hDC98;
defparam \Mux57~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N4
cycloneive_lcell_comb \rfile[31][6]~feeder (
// Equation(s):
// \rfile[31][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[31][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[31][6]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[31][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y31_N5
dffeas \rfile[31][6] (
	.clk(!CLK),
	.d(\rfile[31][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][6] .is_wysiwyg = "true";
defparam \rfile[31][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N23
dffeas \rfile[23][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][6] .is_wysiwyg = "true";
defparam \rfile[23][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y29_N25
dffeas \rfile[27][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][6] .is_wysiwyg = "true";
defparam \rfile[27][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N5
dffeas \rfile[19][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][6] .is_wysiwyg = "true";
defparam \rfile[19][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N24
cycloneive_lcell_comb \Mux57~7 (
// Equation(s):
// \Mux57~7_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[27][6]~q )) # (!instruction_D[19] & ((\rfile[19][6]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[27][6]~q ),
	.datad(\rfile[19][6]~q ),
	.cin(gnd),
	.combout(\Mux57~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~7 .lut_mask = 16'hD9C8;
defparam \Mux57~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N22
cycloneive_lcell_comb \Mux57~8 (
// Equation(s):
// \Mux57~8_combout  = (instruction_D[18] & ((\Mux57~7_combout  & (\rfile[31][6]~q )) # (!\Mux57~7_combout  & ((\rfile[23][6]~q ))))) # (!instruction_D[18] & (((\Mux57~7_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[31][6]~q ),
	.datac(\rfile[23][6]~q ),
	.datad(\Mux57~7_combout ),
	.cin(gnd),
	.combout(\Mux57~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~8 .lut_mask = 16'hDDA0;
defparam \Mux57~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N16
cycloneive_lcell_comb \rfile[7][6]~feeder (
// Equation(s):
// \rfile[7][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_6),
	.cin(gnd),
	.combout(\rfile[7][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[7][6]~feeder .lut_mask = 16'hFF00;
defparam \rfile[7][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y27_N17
dffeas \rfile[7][6] (
	.clk(!CLK),
	.d(\rfile[7][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][6] .is_wysiwyg = "true";
defparam \rfile[7][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N13
dffeas \rfile[5][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][6] .is_wysiwyg = "true";
defparam \rfile[5][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N12
cycloneive_lcell_comb \Mux57~10 (
// Equation(s):
// \Mux57~10_combout  = (instruction_D[16] & (((\rfile[5][6]~q ) # (instruction_D[17])))) # (!instruction_D[16] & (\rfile[4][6]~q  & ((!instruction_D[17]))))

	.dataa(\rfile[4][6]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[5][6]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux57~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~10 .lut_mask = 16'hCCE2;
defparam \Mux57~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N22
cycloneive_lcell_comb \rfile[6][6]~feeder (
// Equation(s):
// \rfile[6][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_6),
	.cin(gnd),
	.combout(\rfile[6][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][6]~feeder .lut_mask = 16'hFF00;
defparam \rfile[6][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y27_N23
dffeas \rfile[6][6] (
	.clk(!CLK),
	.d(\rfile[6][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][6] .is_wysiwyg = "true";
defparam \rfile[6][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N18
cycloneive_lcell_comb \Mux57~11 (
// Equation(s):
// \Mux57~11_combout  = (instruction_D[17] & ((\Mux57~10_combout  & (\rfile[7][6]~q )) # (!\Mux57~10_combout  & ((\rfile[6][6]~q ))))) # (!instruction_D[17] & (((\Mux57~10_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[7][6]~q ),
	.datac(\Mux57~10_combout ),
	.datad(\rfile[6][6]~q ),
	.cin(gnd),
	.combout(\Mux57~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~11 .lut_mask = 16'hDAD0;
defparam \Mux57~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N10
cycloneive_lcell_comb \rfile[14][6]~feeder (
// Equation(s):
// \rfile[14][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[14][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[14][6]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[14][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N11
dffeas \rfile[14][6] (
	.clk(!CLK),
	.d(\rfile[14][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][6] .is_wysiwyg = "true";
defparam \rfile[14][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N31
dffeas \rfile[12][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][6] .is_wysiwyg = "true";
defparam \rfile[12][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N13
dffeas \rfile[13][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][6] .is_wysiwyg = "true";
defparam \rfile[13][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N30
cycloneive_lcell_comb \Mux57~17 (
// Equation(s):
// \Mux57~17_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][6]~q ))) # (!instruction_D[16] & (\rfile[12][6]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[12][6]~q ),
	.datad(\rfile[13][6]~q ),
	.cin(gnd),
	.combout(\Mux57~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~17 .lut_mask = 16'hDC98;
defparam \Mux57~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N28
cycloneive_lcell_comb \rfile[15][6]~feeder (
// Equation(s):
// \rfile[15][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_6),
	.cin(gnd),
	.combout(\rfile[15][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][6]~feeder .lut_mask = 16'hFF00;
defparam \rfile[15][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N29
dffeas \rfile[15][6] (
	.clk(!CLK),
	.d(\rfile[15][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][6] .is_wysiwyg = "true";
defparam \rfile[15][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N18
cycloneive_lcell_comb \Mux57~18 (
// Equation(s):
// \Mux57~18_combout  = (instruction_D[17] & ((\Mux57~17_combout  & ((\rfile[15][6]~q ))) # (!\Mux57~17_combout  & (\rfile[14][6]~q )))) # (!instruction_D[17] & (((\Mux57~17_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[14][6]~q ),
	.datac(\Mux57~17_combout ),
	.datad(\rfile[15][6]~q ),
	.cin(gnd),
	.combout(\Mux57~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~18 .lut_mask = 16'hF858;
defparam \Mux57~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N6
cycloneive_lcell_comb \rfile[2][6]~feeder (
// Equation(s):
// \rfile[2][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_6),
	.cin(gnd),
	.combout(\rfile[2][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][6]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y27_N7
dffeas \rfile[2][6] (
	.clk(!CLK),
	.d(\rfile[2][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][6] .is_wysiwyg = "true";
defparam \rfile[2][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N14
cycloneive_lcell_comb \rfile[1][6]~feeder (
// Equation(s):
// \rfile[1][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[1][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[1][6]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[1][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N15
dffeas \rfile[1][6] (
	.clk(!CLK),
	.d(\rfile[1][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][6] .is_wysiwyg = "true";
defparam \rfile[1][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N20
cycloneive_lcell_comb \rfile[3][6]~feeder (
// Equation(s):
// \rfile[3][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[3][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[3][6]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[3][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N21
dffeas \rfile[3][6] (
	.clk(!CLK),
	.d(\rfile[3][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][6] .is_wysiwyg = "true";
defparam \rfile[3][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N28
cycloneive_lcell_comb \Mux57~14 (
// Equation(s):
// \Mux57~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][6]~q ))) # (!instruction_D[17] & (\rfile[1][6]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[1][6]~q ),
	.datad(\rfile[3][6]~q ),
	.cin(gnd),
	.combout(\Mux57~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~14 .lut_mask = 16'hA820;
defparam \Mux57~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N22
cycloneive_lcell_comb \Mux57~15 (
// Equation(s):
// \Mux57~15_combout  = (\Mux57~14_combout ) # ((!instruction_D[16] & (instruction_D[17] & \rfile[2][6]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[2][6]~q ),
	.datad(\Mux57~14_combout ),
	.cin(gnd),
	.combout(\Mux57~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~15 .lut_mask = 16'hFF40;
defparam \Mux57~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N27
dffeas \rfile[9][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][6] .is_wysiwyg = "true";
defparam \rfile[9][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N31
dffeas \rfile[10][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][6] .is_wysiwyg = "true";
defparam \rfile[10][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N29
dffeas \rfile[8][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][6] .is_wysiwyg = "true";
defparam \rfile[8][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N30
cycloneive_lcell_comb \Mux57~12 (
// Equation(s):
// \Mux57~12_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\rfile[10][6]~q )) # (!instruction_D[17] & ((\rfile[8][6]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[10][6]~q ),
	.datad(\rfile[8][6]~q ),
	.cin(gnd),
	.combout(\Mux57~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~12 .lut_mask = 16'hD9C8;
defparam \Mux57~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N26
cycloneive_lcell_comb \Mux57~13 (
// Equation(s):
// \Mux57~13_combout  = (instruction_D[16] & ((\Mux57~12_combout  & (\rfile[11][6]~q )) # (!\Mux57~12_combout  & ((\rfile[9][6]~q ))))) # (!instruction_D[16] & (((\Mux57~12_combout ))))

	.dataa(\rfile[11][6]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[9][6]~q ),
	.datad(\Mux57~12_combout ),
	.cin(gnd),
	.combout(\Mux57~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~13 .lut_mask = 16'hBBC0;
defparam \Mux57~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N0
cycloneive_lcell_comb \Mux57~16 (
// Equation(s):
// \Mux57~16_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\Mux57~13_combout )))) # (!instruction_D[19] & (!instruction_D[18] & (\Mux57~15_combout )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux57~15_combout ),
	.datad(\Mux57~13_combout ),
	.cin(gnd),
	.combout(\Mux57~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~16 .lut_mask = 16'hBA98;
defparam \Mux57~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y27_N2
cycloneive_lcell_comb \rfile[27][5]~feeder (
// Equation(s):
// \rfile[27][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_5),
	.cin(gnd),
	.combout(\rfile[27][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[27][5]~feeder .lut_mask = 16'hFF00;
defparam \rfile[27][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y27_N3
dffeas \rfile[27][5] (
	.clk(!CLK),
	.d(\rfile[27][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][5] .is_wysiwyg = "true";
defparam \rfile[27][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y27_N18
cycloneive_lcell_comb \rfile[19][5]~feeder (
// Equation(s):
// \rfile[19][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_5),
	.cin(gnd),
	.combout(\rfile[19][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[19][5]~feeder .lut_mask = 16'hFF00;
defparam \rfile[19][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y27_N19
dffeas \rfile[19][5] (
	.clk(!CLK),
	.d(\rfile[19][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][5] .is_wysiwyg = "true";
defparam \rfile[19][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y27_N0
cycloneive_lcell_comb \rfile[23][5]~feeder (
// Equation(s):
// \rfile[23][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_5),
	.cin(gnd),
	.combout(\rfile[23][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[23][5]~feeder .lut_mask = 16'hFF00;
defparam \rfile[23][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y27_N1
dffeas \rfile[23][5] (
	.clk(!CLK),
	.d(\rfile[23][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][5] .is_wysiwyg = "true";
defparam \rfile[23][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y27_N12
cycloneive_lcell_comb \Mux58~7 (
// Equation(s):
// \Mux58~7_combout  = (instruction_D[18] & (((instruction_D[19]) # (\rfile[23][5]~q )))) # (!instruction_D[18] & (\rfile[19][5]~q  & (!instruction_D[19])))

	.dataa(instruction_D_18),
	.datab(\rfile[19][5]~q ),
	.datac(instruction_D_19),
	.datad(\rfile[23][5]~q ),
	.cin(gnd),
	.combout(\Mux58~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~7 .lut_mask = 16'hAEA4;
defparam \Mux58~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N18
cycloneive_lcell_comb \rfile[31][5]~feeder (
// Equation(s):
// \rfile[31][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_5),
	.cin(gnd),
	.combout(\rfile[31][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[31][5]~feeder .lut_mask = 16'hFF00;
defparam \rfile[31][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y31_N19
dffeas \rfile[31][5] (
	.clk(!CLK),
	.d(\rfile[31][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][5] .is_wysiwyg = "true";
defparam \rfile[31][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y27_N12
cycloneive_lcell_comb \Mux58~8 (
// Equation(s):
// \Mux58~8_combout  = (instruction_D[19] & ((\Mux58~7_combout  & ((\rfile[31][5]~q ))) # (!\Mux58~7_combout  & (\rfile[27][5]~q )))) # (!instruction_D[19] & (((\Mux58~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[27][5]~q ),
	.datac(\Mux58~7_combout ),
	.datad(\rfile[31][5]~q ),
	.cin(gnd),
	.combout(\Mux58~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~8 .lut_mask = 16'hF858;
defparam \Mux58~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y28_N11
dffeas \rfile[17][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][5] .is_wysiwyg = "true";
defparam \rfile[17][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N3
dffeas \rfile[21][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][5] .is_wysiwyg = "true";
defparam \rfile[21][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N10
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[21][5]~q ))) # (!instruction_D[18] & (\rfile[17][5]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[17][5]~q ),
	.datad(\rfile[21][5]~q ),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'hDC98;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N21
dffeas \rfile[29][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][5] .is_wysiwyg = "true";
defparam \rfile[29][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N13
dffeas \rfile[25][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][5] .is_wysiwyg = "true";
defparam \rfile[25][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N12
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (\Mux58~0_combout  & ((\rfile[29][5]~q ) # ((!instruction_D[19])))) # (!\Mux58~0_combout  & (((\rfile[25][5]~q  & instruction_D[19]))))

	.dataa(\Mux58~0_combout ),
	.datab(\rfile[29][5]~q ),
	.datac(\rfile[25][5]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hD8AA;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y32_N3
dffeas \rfile[20][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][5] .is_wysiwyg = "true";
defparam \rfile[20][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N13
dffeas \rfile[24][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][5] .is_wysiwyg = "true";
defparam \rfile[24][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N3
dffeas \rfile[16][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][5] .is_wysiwyg = "true";
defparam \rfile[16][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N12
cycloneive_lcell_comb \Mux58~4 (
// Equation(s):
// \Mux58~4_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[24][5]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[16][5]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[24][5]~q ),
	.datad(\rfile[16][5]~q ),
	.cin(gnd),
	.combout(\Mux58~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~4 .lut_mask = 16'hB9A8;
defparam \Mux58~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N2
cycloneive_lcell_comb \Mux58~5 (
// Equation(s):
// \Mux58~5_combout  = (instruction_D[18] & ((\Mux58~4_combout  & (\rfile[28][5]~q )) # (!\Mux58~4_combout  & ((\rfile[20][5]~q ))))) # (!instruction_D[18] & (((\Mux58~4_combout ))))

	.dataa(\rfile[28][5]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[20][5]~q ),
	.datad(\Mux58~4_combout ),
	.cin(gnd),
	.combout(\Mux58~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~5 .lut_mask = 16'hBBC0;
defparam \Mux58~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y36_N25
dffeas \rfile[30][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][5] .is_wysiwyg = "true";
defparam \rfile[30][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y36_N19
dffeas \rfile[26][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][5] .is_wysiwyg = "true";
defparam \rfile[26][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N18
cycloneive_lcell_comb \Mux58~2 (
// Equation(s):
// \Mux58~2_combout  = (instruction_D[19] & (((\rfile[26][5]~q ) # (instruction_D[18])))) # (!instruction_D[19] & (\rfile[18][5]~q  & ((!instruction_D[18]))))

	.dataa(\rfile[18][5]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[26][5]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux58~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~2 .lut_mask = 16'hCCE2;
defparam \Mux58~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N24
cycloneive_lcell_comb \Mux58~3 (
// Equation(s):
// \Mux58~3_combout  = (instruction_D[18] & ((\Mux58~2_combout  & ((\rfile[30][5]~q ))) # (!\Mux58~2_combout  & (\rfile[22][5]~q )))) # (!instruction_D[18] & (((\Mux58~2_combout ))))

	.dataa(\rfile[22][5]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[30][5]~q ),
	.datad(\Mux58~2_combout ),
	.cin(gnd),
	.combout(\Mux58~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~3 .lut_mask = 16'hF388;
defparam \Mux58~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N18
cycloneive_lcell_comb \Mux58~6 (
// Equation(s):
// \Mux58~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux58~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & (\Mux58~5_combout )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux58~5_combout ),
	.datad(\Mux58~3_combout ),
	.cin(gnd),
	.combout(\Mux58~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~6 .lut_mask = 16'hBA98;
defparam \Mux58~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N28
cycloneive_lcell_comb \rfile[11][5]~feeder (
// Equation(s):
// \rfile[11][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[11][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][5]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[11][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y27_N29
dffeas \rfile[11][5] (
	.clk(!CLK),
	.d(\rfile[11][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][5] .is_wysiwyg = "true";
defparam \rfile[11][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N11
dffeas \rfile[10][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][5] .is_wysiwyg = "true";
defparam \rfile[10][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N13
dffeas \rfile[8][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][5] .is_wysiwyg = "true";
defparam \rfile[8][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N10
cycloneive_lcell_comb \Mux58~10 (
// Equation(s):
// \Mux58~10_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\rfile[10][5]~q )) # (!instruction_D[17] & ((\rfile[8][5]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[10][5]~q ),
	.datad(\rfile[8][5]~q ),
	.cin(gnd),
	.combout(\Mux58~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~10 .lut_mask = 16'hD9C8;
defparam \Mux58~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N24
cycloneive_lcell_comb \rfile[9][5]~feeder (
// Equation(s):
// \rfile[9][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_5),
	.cin(gnd),
	.combout(\rfile[9][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][5]~feeder .lut_mask = 16'hFF00;
defparam \rfile[9][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N25
dffeas \rfile[9][5] (
	.clk(!CLK),
	.d(\rfile[9][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][5] .is_wysiwyg = "true";
defparam \rfile[9][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N22
cycloneive_lcell_comb \Mux58~11 (
// Equation(s):
// \Mux58~11_combout  = (instruction_D[16] & ((\Mux58~10_combout  & (\rfile[11][5]~q )) # (!\Mux58~10_combout  & ((\rfile[9][5]~q ))))) # (!instruction_D[16] & (((\Mux58~10_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][5]~q ),
	.datac(\Mux58~10_combout ),
	.datad(\rfile[9][5]~q ),
	.cin(gnd),
	.combout(\Mux58~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~11 .lut_mask = 16'hDAD0;
defparam \Mux58~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N4
cycloneive_lcell_comb \rfile[15][5]~feeder (
// Equation(s):
// \rfile[15][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[15][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][5]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[15][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N5
dffeas \rfile[15][5] (
	.clk(!CLK),
	.d(\rfile[15][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][5] .is_wysiwyg = "true";
defparam \rfile[15][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N21
dffeas \rfile[14][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][5] .is_wysiwyg = "true";
defparam \rfile[14][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N7
dffeas \rfile[13][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][5] .is_wysiwyg = "true";
defparam \rfile[13][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N1
dffeas \rfile[12][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][5] .is_wysiwyg = "true";
defparam \rfile[12][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N6
cycloneive_lcell_comb \Mux58~17 (
// Equation(s):
// \Mux58~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][5]~q )))) # (!instruction_D[16] & (!instruction_D[17] & ((\rfile[12][5]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[13][5]~q ),
	.datad(\rfile[12][5]~q ),
	.cin(gnd),
	.combout(\Mux58~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~17 .lut_mask = 16'hB9A8;
defparam \Mux58~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N20
cycloneive_lcell_comb \Mux58~18 (
// Equation(s):
// \Mux58~18_combout  = (instruction_D[17] & ((\Mux58~17_combout  & (\rfile[15][5]~q )) # (!\Mux58~17_combout  & ((\rfile[14][5]~q ))))) # (!instruction_D[17] & (((\Mux58~17_combout ))))

	.dataa(\rfile[15][5]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[14][5]~q ),
	.datad(\Mux58~17_combout ),
	.cin(gnd),
	.combout(\Mux58~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~18 .lut_mask = 16'hBBC0;
defparam \Mux58~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N26
cycloneive_lcell_comb \rfile[3][5]~feeder (
// Equation(s):
// \rfile[3][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_5),
	.cin(gnd),
	.combout(\rfile[3][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[3][5]~feeder .lut_mask = 16'hFF00;
defparam \rfile[3][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N27
dffeas \rfile[3][5] (
	.clk(!CLK),
	.d(\rfile[3][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][5] .is_wysiwyg = "true";
defparam \rfile[3][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N12
cycloneive_lcell_comb \rfile[1][5]~feeder (
// Equation(s):
// \rfile[1][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_5),
	.cin(gnd),
	.combout(\rfile[1][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[1][5]~feeder .lut_mask = 16'hFF00;
defparam \rfile[1][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N13
dffeas \rfile[1][5] (
	.clk(!CLK),
	.d(\rfile[1][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][5] .is_wysiwyg = "true";
defparam \rfile[1][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N10
cycloneive_lcell_comb \Mux58~14 (
// Equation(s):
// \Mux58~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][5]~q )) # (!instruction_D[17] & ((\rfile[1][5]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[3][5]~q ),
	.datad(\rfile[1][5]~q ),
	.cin(gnd),
	.combout(\Mux58~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~14 .lut_mask = 16'hC480;
defparam \Mux58~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N24
cycloneive_lcell_comb \rfile[2][5]~feeder (
// Equation(s):
// \rfile[2][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[2][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][5]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[2][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y27_N25
dffeas \rfile[2][5] (
	.clk(!CLK),
	.d(\rfile[2][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][5] .is_wysiwyg = "true";
defparam \rfile[2][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N14
cycloneive_lcell_comb \Mux58~15 (
// Equation(s):
// \Mux58~15_combout  = (\Mux58~14_combout ) # ((!instruction_D[16] & (instruction_D[17] & \rfile[2][5]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux58~14_combout ),
	.datad(\rfile[2][5]~q ),
	.cin(gnd),
	.combout(\Mux58~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~15 .lut_mask = 16'hF4F0;
defparam \Mux58~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N8
cycloneive_lcell_comb \rfile[6][5]~feeder (
// Equation(s):
// \rfile[6][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_5),
	.cin(gnd),
	.combout(\rfile[6][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][5]~feeder .lut_mask = 16'hFF00;
defparam \rfile[6][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y27_N9
dffeas \rfile[6][5] (
	.clk(!CLK),
	.d(\rfile[6][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][5] .is_wysiwyg = "true";
defparam \rfile[6][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N14
cycloneive_lcell_comb \rfile[7][5]~feeder (
// Equation(s):
// \rfile[7][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_5),
	.cin(gnd),
	.combout(\rfile[7][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[7][5]~feeder .lut_mask = 16'hFF00;
defparam \rfile[7][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y27_N15
dffeas \rfile[7][5] (
	.clk(!CLK),
	.d(\rfile[7][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][5] .is_wysiwyg = "true";
defparam \rfile[7][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N25
dffeas \rfile[5][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][5] .is_wysiwyg = "true";
defparam \rfile[5][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N19
dffeas \rfile[4][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][5] .is_wysiwyg = "true";
defparam \rfile[4][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N24
cycloneive_lcell_comb \Mux58~12 (
// Equation(s):
// \Mux58~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[5][5]~q )) # (!instruction_D[16] & ((\rfile[4][5]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[5][5]~q ),
	.datad(\rfile[4][5]~q ),
	.cin(gnd),
	.combout(\Mux58~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~12 .lut_mask = 16'hD9C8;
defparam \Mux58~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N28
cycloneive_lcell_comb \Mux58~13 (
// Equation(s):
// \Mux58~13_combout  = (instruction_D[17] & ((\Mux58~12_combout  & ((\rfile[7][5]~q ))) # (!\Mux58~12_combout  & (\rfile[6][5]~q )))) # (!instruction_D[17] & (((\Mux58~12_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[6][5]~q ),
	.datac(\rfile[7][5]~q ),
	.datad(\Mux58~12_combout ),
	.cin(gnd),
	.combout(\Mux58~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~13 .lut_mask = 16'hF588;
defparam \Mux58~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N12
cycloneive_lcell_comb \Mux58~16 (
// Equation(s):
// \Mux58~16_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\Mux58~13_combout )))) # (!instruction_D[18] & (!instruction_D[19] & (\Mux58~15_combout )))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\Mux58~15_combout ),
	.datad(\Mux58~13_combout ),
	.cin(gnd),
	.combout(\Mux58~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~16 .lut_mask = 16'hBA98;
defparam \Mux58~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N23
dffeas \rfile[21][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][2] .is_wysiwyg = "true";
defparam \rfile[21][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N18
cycloneive_lcell_comb \rfile[17][2]~feeder (
// Equation(s):
// \rfile[17][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[17][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[17][2]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[17][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y28_N19
dffeas \rfile[17][2] (
	.clk(!CLK),
	.d(\rfile[17][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][2] .is_wysiwyg = "true";
defparam \rfile[17][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N22
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[21][2]~q )) # (!instruction_D[23] & ((\rfile[17][2]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[21][2]~q ),
	.datad(\rfile[17][2]~q ),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hD9C8;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N5
dffeas \rfile[29][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][2] .is_wysiwyg = "true";
defparam \rfile[29][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N21
dffeas \rfile[25][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][2] .is_wysiwyg = "true";
defparam \rfile[25][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N4
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (\Mux29~0_combout  & (((\rfile[29][2]~q )) # (!instruction_D[24]))) # (!\Mux29~0_combout  & (instruction_D[24] & ((\rfile[25][2]~q ))))

	.dataa(\Mux29~0_combout ),
	.datab(instruction_D_24),
	.datac(\rfile[29][2]~q ),
	.datad(\rfile[25][2]~q ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hE6A2;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N14
cycloneive_lcell_comb \rfile[23][2]~feeder (
// Equation(s):
// \rfile[23][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[23][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[23][2]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[23][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y29_N15
dffeas \rfile[23][2] (
	.clk(!CLK),
	.d(\rfile[23][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][2] .is_wysiwyg = "true";
defparam \rfile[23][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y29_N27
dffeas \rfile[19][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][2] .is_wysiwyg = "true";
defparam \rfile[19][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N28
cycloneive_lcell_comb \Mux29~7 (
// Equation(s):
// \Mux29~7_combout  = (instruction_D[24] & (((instruction_D[23])))) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[23][2]~q )) # (!instruction_D[23] & ((\rfile[19][2]~q )))))

	.dataa(instruction_D_24),
	.datab(\rfile[23][2]~q ),
	.datac(instruction_D_23),
	.datad(\rfile[19][2]~q ),
	.cin(gnd),
	.combout(\Mux29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~7 .lut_mask = 16'hE5E0;
defparam \Mux29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y29_N3
dffeas \rfile[31][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][2] .is_wysiwyg = "true";
defparam \rfile[31][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y29_N7
dffeas \rfile[27][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][2] .is_wysiwyg = "true";
defparam \rfile[27][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N2
cycloneive_lcell_comb \Mux29~8 (
// Equation(s):
// \Mux29~8_combout  = (instruction_D[24] & ((\Mux29~7_combout  & (\rfile[31][2]~q )) # (!\Mux29~7_combout  & ((\rfile[27][2]~q ))))) # (!instruction_D[24] & (\Mux29~7_combout ))

	.dataa(instruction_D_24),
	.datab(\Mux29~7_combout ),
	.datac(\rfile[31][2]~q ),
	.datad(\rfile[27][2]~q ),
	.cin(gnd),
	.combout(\Mux29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~8 .lut_mask = 16'hE6C4;
defparam \Mux29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y36_N25
dffeas \rfile[30][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][2] .is_wysiwyg = "true";
defparam \rfile[30][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y36_N10
cycloneive_lcell_comb \rfile[22][2]~feeder (
// Equation(s):
// \rfile[22][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_2),
	.cin(gnd),
	.combout(\rfile[22][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[22][2]~feeder .lut_mask = 16'hFF00;
defparam \rfile[22][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y36_N11
dffeas \rfile[22][2] (
	.clk(!CLK),
	.d(\rfile[22][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][2] .is_wysiwyg = "true";
defparam \rfile[22][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y36_N8
cycloneive_lcell_comb \rfile[18][2]~feeder (
// Equation(s):
// \rfile[18][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_2),
	.cin(gnd),
	.combout(\rfile[18][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[18][2]~feeder .lut_mask = 16'hFF00;
defparam \rfile[18][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y36_N9
dffeas \rfile[18][2] (
	.clk(!CLK),
	.d(\rfile[18][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][2] .is_wysiwyg = "true";
defparam \rfile[18][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N20
cycloneive_lcell_comb \rfile[26][2]~feeder (
// Equation(s):
// \rfile[26][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[26][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[26][2]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[26][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y36_N21
dffeas \rfile[26][2] (
	.clk(!CLK),
	.d(\rfile[26][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][2] .is_wysiwyg = "true";
defparam \rfile[26][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N10
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][2]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[18][2]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][2]~q ),
	.datad(\rfile[26][2]~q ),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hBA98;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N26
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (instruction_D[23] & ((\Mux29~2_combout  & (\rfile[30][2]~q )) # (!\Mux29~2_combout  & ((\rfile[22][2]~q ))))) # (!instruction_D[23] & (((\Mux29~2_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[30][2]~q ),
	.datac(\rfile[22][2]~q ),
	.datad(\Mux29~2_combout ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'hDDA0;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y32_N9
dffeas \rfile[20][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][2] .is_wysiwyg = "true";
defparam \rfile[20][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N6
cycloneive_lcell_comb \rfile[16][2]~feeder (
// Equation(s):
// \rfile[16][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[16][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[16][2]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[16][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y32_N7
dffeas \rfile[16][2] (
	.clk(!CLK),
	.d(\rfile[16][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][2] .is_wysiwyg = "true";
defparam \rfile[16][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X77_Y32_N18
cycloneive_lcell_comb \rfile[24][2]~feeder (
// Equation(s):
// \rfile[24][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_2),
	.cin(gnd),
	.combout(\rfile[24][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[24][2]~feeder .lut_mask = 16'hFF00;
defparam \rfile[24][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X77_Y32_N19
dffeas \rfile[24][2] (
	.clk(!CLK),
	.d(\rfile[24][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][2] .is_wysiwyg = "true";
defparam \rfile[24][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X77_Y32_N24
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[24][2]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[16][2]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[16][2]~q ),
	.datad(\rfile[24][2]~q ),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'hBA98;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y32_N12
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (instruction_D[23] & ((\Mux29~4_combout  & (\rfile[28][2]~q )) # (!\Mux29~4_combout  & ((\rfile[20][2]~q ))))) # (!instruction_D[23] & (((\Mux29~4_combout ))))

	.dataa(\rfile[28][2]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[20][2]~q ),
	.datad(\Mux29~4_combout ),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'hBBC0;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N24
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// \Mux29~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\Mux29~3_combout )) # (!instruction_D[22] & ((\Mux29~5_combout )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux29~3_combout ),
	.datad(\Mux29~5_combout ),
	.cin(gnd),
	.combout(\Mux29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hD9C8;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N14
cycloneive_lcell_comb \rfile[9][2]~feeder (
// Equation(s):
// \rfile[9][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_2),
	.cin(gnd),
	.combout(\rfile[9][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][2]~feeder .lut_mask = 16'hFF00;
defparam \rfile[9][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N15
dffeas \rfile[9][2] (
	.clk(!CLK),
	.d(\rfile[9][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][2] .is_wysiwyg = "true";
defparam \rfile[9][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N4
cycloneive_lcell_comb \rfile[11][2]~feeder (
// Equation(s):
// \rfile[11][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_2),
	.cin(gnd),
	.combout(\rfile[11][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][2]~feeder .lut_mask = 16'hFF00;
defparam \rfile[11][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N5
dffeas \rfile[11][2] (
	.clk(!CLK),
	.d(\rfile[11][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][2] .is_wysiwyg = "true";
defparam \rfile[11][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N27
dffeas \rfile[10][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][2] .is_wysiwyg = "true";
defparam \rfile[10][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N6
cycloneive_lcell_comb \rfile[8][2]~feeder (
// Equation(s):
// \rfile[8][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_2),
	.cin(gnd),
	.combout(\rfile[8][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[8][2]~feeder .lut_mask = 16'hFF00;
defparam \rfile[8][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N7
dffeas \rfile[8][2] (
	.clk(!CLK),
	.d(\rfile[8][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][2] .is_wysiwyg = "true";
defparam \rfile[8][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N26
cycloneive_lcell_comb \Mux29~10 (
// Equation(s):
// \Mux29~10_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][2]~q )))) # (!instruction_D[22] & (!instruction_D[21] & ((\rfile[8][2]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[10][2]~q ),
	.datad(\rfile[8][2]~q ),
	.cin(gnd),
	.combout(\Mux29~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~10 .lut_mask = 16'hB9A8;
defparam \Mux29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N2
cycloneive_lcell_comb \Mux29~11 (
// Equation(s):
// \Mux29~11_combout  = (instruction_D[21] & ((\Mux29~10_combout  & ((\rfile[11][2]~q ))) # (!\Mux29~10_combout  & (\rfile[9][2]~q )))) # (!instruction_D[21] & (((\Mux29~10_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[9][2]~q ),
	.datac(\rfile[11][2]~q ),
	.datad(\Mux29~10_combout ),
	.cin(gnd),
	.combout(\Mux29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~11 .lut_mask = 16'hF588;
defparam \Mux29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N14
cycloneive_lcell_comb \rfile[15][2]~feeder (
// Equation(s):
// \rfile[15][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_2),
	.cin(gnd),
	.combout(\rfile[15][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][2]~feeder .lut_mask = 16'hFF00;
defparam \rfile[15][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N15
dffeas \rfile[15][2] (
	.clk(!CLK),
	.d(\rfile[15][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][2] .is_wysiwyg = "true";
defparam \rfile[15][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N1
dffeas \rfile[14][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][2] .is_wysiwyg = "true";
defparam \rfile[14][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N30
cycloneive_lcell_comb \rfile[13][2]~feeder (
// Equation(s):
// \rfile[13][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[13][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[13][2]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[13][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N31
dffeas \rfile[13][2] (
	.clk(!CLK),
	.d(\rfile[13][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][2] .is_wysiwyg = "true";
defparam \rfile[13][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N13
dffeas \rfile[12][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][2] .is_wysiwyg = "true";
defparam \rfile[12][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N12
cycloneive_lcell_comb \Mux29~17 (
// Equation(s):
// \Mux29~17_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][2]~q )) # (!instruction_D[21] & ((\rfile[12][2]~q )))))

	.dataa(instruction_D_22),
	.datab(\rfile[13][2]~q ),
	.datac(\rfile[12][2]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux29~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~17 .lut_mask = 16'hEE50;
defparam \Mux29~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N26
cycloneive_lcell_comb \Mux29~18 (
// Equation(s):
// \Mux29~18_combout  = (instruction_D[22] & ((\Mux29~17_combout  & (\rfile[15][2]~q )) # (!\Mux29~17_combout  & ((\rfile[14][2]~q ))))) # (!instruction_D[22] & (((\Mux29~17_combout ))))

	.dataa(\rfile[15][2]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[14][2]~q ),
	.datad(\Mux29~17_combout ),
	.cin(gnd),
	.combout(\Mux29~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~18 .lut_mask = 16'hBBC0;
defparam \Mux29~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N17
dffeas \rfile[6][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][2] .is_wysiwyg = "true";
defparam \rfile[6][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N23
dffeas \rfile[7][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][2] .is_wysiwyg = "true";
defparam \rfile[7][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N29
dffeas \rfile[5][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][2] .is_wysiwyg = "true";
defparam \rfile[5][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N11
dffeas \rfile[4][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][2] .is_wysiwyg = "true";
defparam \rfile[4][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N28
cycloneive_lcell_comb \Mux29~12 (
// Equation(s):
// \Mux29~12_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[5][2]~q )) # (!instruction_D[21] & ((\rfile[4][2]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[5][2]~q ),
	.datad(\rfile[4][2]~q ),
	.cin(gnd),
	.combout(\Mux29~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~12 .lut_mask = 16'hD9C8;
defparam \Mux29~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N22
cycloneive_lcell_comb \Mux29~13 (
// Equation(s):
// \Mux29~13_combout  = (instruction_D[22] & ((\Mux29~12_combout  & ((\rfile[7][2]~q ))) # (!\Mux29~12_combout  & (\rfile[6][2]~q )))) # (!instruction_D[22] & (((\Mux29~12_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[6][2]~q ),
	.datac(\rfile[7][2]~q ),
	.datad(\Mux29~12_combout ),
	.cin(gnd),
	.combout(\Mux29~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~13 .lut_mask = 16'hF588;
defparam \Mux29~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N16
cycloneive_lcell_comb \rfile[2][2]~feeder (
// Equation(s):
// \rfile[2][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_2),
	.cin(gnd),
	.combout(\rfile[2][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][2]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N17
dffeas \rfile[2][2] (
	.clk(!CLK),
	.d(\rfile[2][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][2] .is_wysiwyg = "true";
defparam \rfile[2][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N15
dffeas \rfile[1][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][2] .is_wysiwyg = "true";
defparam \rfile[1][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N12
cycloneive_lcell_comb \rfile[3][2]~feeder (
// Equation(s):
// \rfile[3][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[3][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[3][2]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[3][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N13
dffeas \rfile[3][2] (
	.clk(!CLK),
	.d(\rfile[3][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][2] .is_wysiwyg = "true";
defparam \rfile[3][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N20
cycloneive_lcell_comb \Mux29~14 (
// Equation(s):
// \Mux29~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][2]~q ))) # (!instruction_D[22] & (\rfile[1][2]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[1][2]~q ),
	.datad(\rfile[3][2]~q ),
	.cin(gnd),
	.combout(\Mux29~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~14 .lut_mask = 16'hA820;
defparam \Mux29~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N22
cycloneive_lcell_comb \Mux29~15 (
// Equation(s):
// \Mux29~15_combout  = (\Mux29~14_combout ) # ((!instruction_D[21] & (\rfile[2][2]~q  & instruction_D[22])))

	.dataa(instruction_D_21),
	.datab(\rfile[2][2]~q ),
	.datac(instruction_D_22),
	.datad(\Mux29~14_combout ),
	.cin(gnd),
	.combout(\Mux29~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~15 .lut_mask = 16'hFF40;
defparam \Mux29~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N12
cycloneive_lcell_comb \Mux29~16 (
// Equation(s):
// \Mux29~16_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\Mux29~13_combout )))) # (!instruction_D[23] & (!instruction_D[24] & ((\Mux29~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux29~13_combout ),
	.datad(\Mux29~15_combout ),
	.cin(gnd),
	.combout(\Mux29~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~16 .lut_mask = 16'hB9A8;
defparam \Mux29~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y33_N25
dffeas \rfile[16][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][1] .is_wysiwyg = "true";
defparam \rfile[16][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y33_N27
dffeas \rfile[24][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][1] .is_wysiwyg = "true";
defparam \rfile[24][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N24
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// \Mux30~4_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\rfile[24][1]~q ))) # (!instruction_D[24] & (\rfile[16][1]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[16][1]~q ),
	.datad(\rfile[24][1]~q ),
	.cin(gnd),
	.combout(\Mux30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'hDC98;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N25
dffeas \rfile[20][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][1] .is_wysiwyg = "true";
defparam \rfile[20][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N2
cycloneive_lcell_comb \rfile[28][1]~feeder (
// Equation(s):
// \rfile[28][1]~feeder_combout  = \wdat_WB[1]~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[28][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][1]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[28][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N3
dffeas \rfile[28][1] (
	.clk(!CLK),
	.d(\rfile[28][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][1] .is_wysiwyg = "true";
defparam \rfile[28][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N24
cycloneive_lcell_comb \Mux30~5 (
// Equation(s):
// \Mux30~5_combout  = (instruction_D[23] & ((\Mux30~4_combout  & ((\rfile[28][1]~q ))) # (!\Mux30~4_combout  & (\rfile[20][1]~q )))) # (!instruction_D[23] & (\Mux30~4_combout ))

	.dataa(instruction_D_23),
	.datab(\Mux30~4_combout ),
	.datac(\rfile[20][1]~q ),
	.datad(\rfile[28][1]~q ),
	.cin(gnd),
	.combout(\Mux30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~5 .lut_mask = 16'hEC64;
defparam \Mux30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y35_N15
dffeas \rfile[22][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][1] .is_wysiwyg = "true";
defparam \rfile[22][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y35_N25
dffeas \rfile[30][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][1] .is_wysiwyg = "true";
defparam \rfile[30][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N14
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (\Mux30~2_combout  & (((\rfile[30][1]~q )) # (!instruction_D[23]))) # (!\Mux30~2_combout  & (instruction_D[23] & (\rfile[22][1]~q )))

	.dataa(\Mux30~2_combout ),
	.datab(instruction_D_23),
	.datac(\rfile[22][1]~q ),
	.datad(\rfile[30][1]~q ),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'hEA62;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N16
cycloneive_lcell_comb \Mux30~6 (
// Equation(s):
// \Mux30~6_combout  = (instruction_D[21] & (((instruction_D[22])))) # (!instruction_D[21] & ((instruction_D[22] & ((\Mux30~3_combout ))) # (!instruction_D[22] & (\Mux30~5_combout ))))

	.dataa(instruction_D_21),
	.datab(\Mux30~5_combout ),
	.datac(instruction_D_22),
	.datad(\Mux30~3_combout ),
	.cin(gnd),
	.combout(\Mux30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~6 .lut_mask = 16'hF4A4;
defparam \Mux30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N9
dffeas \rfile[27][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][1] .is_wysiwyg = "true";
defparam \rfile[27][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y29_N3
dffeas \rfile[31][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][1] .is_wysiwyg = "true";
defparam \rfile[31][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N14
cycloneive_lcell_comb \rfile[23][1]~feeder (
// Equation(s):
// \rfile[23][1]~feeder_combout  = \wdat_WB[1]~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[23][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[23][1]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[23][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N15
dffeas \rfile[23][1] (
	.clk(!CLK),
	.d(\rfile[23][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][1] .is_wysiwyg = "true";
defparam \rfile[23][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N12
cycloneive_lcell_comb \rfile[19][1]~feeder (
// Equation(s):
// \rfile[19][1]~feeder_combout  = \wdat_WB[1]~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[19][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[19][1]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[19][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N13
dffeas \rfile[19][1] (
	.clk(!CLK),
	.d(\rfile[19][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][1] .is_wysiwyg = "true";
defparam \rfile[19][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N22
cycloneive_lcell_comb \Mux30~7 (
// Equation(s):
// \Mux30~7_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[23][1]~q )))) # (!instruction_D[23] & (!instruction_D[24] & ((\rfile[19][1]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[23][1]~q ),
	.datad(\rfile[19][1]~q ),
	.cin(gnd),
	.combout(\Mux30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~7 .lut_mask = 16'hB9A8;
defparam \Mux30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N2
cycloneive_lcell_comb \Mux30~8 (
// Equation(s):
// \Mux30~8_combout  = (instruction_D[24] & ((\Mux30~7_combout  & ((\rfile[31][1]~q ))) # (!\Mux30~7_combout  & (\rfile[27][1]~q )))) # (!instruction_D[24] & (((\Mux30~7_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[27][1]~q ),
	.datac(\rfile[31][1]~q ),
	.datad(\Mux30~7_combout ),
	.cin(gnd),
	.combout(\Mux30~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~8 .lut_mask = 16'hF588;
defparam \Mux30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N1
dffeas \rfile[25][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][1] .is_wysiwyg = "true";
defparam \rfile[25][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N3
dffeas \rfile[29][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][1] .is_wysiwyg = "true";
defparam \rfile[29][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y30_N17
dffeas \rfile[17][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][1] .is_wysiwyg = "true";
defparam \rfile[17][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N16
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (instruction_D[23] & ((\rfile[21][1]~q ) # ((instruction_D[24])))) # (!instruction_D[23] & (((\rfile[17][1]~q  & !instruction_D[24]))))

	.dataa(\rfile[21][1]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[17][1]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hCCB8;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N2
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (instruction_D[24] & ((\Mux30~0_combout  & ((\rfile[29][1]~q ))) # (!\Mux30~0_combout  & (\rfile[25][1]~q )))) # (!instruction_D[24] & (((\Mux30~0_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[25][1]~q ),
	.datac(\rfile[29][1]~q ),
	.datad(\Mux30~0_combout ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hF588;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N13
dffeas \rfile[11][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][1] .is_wysiwyg = "true";
defparam \rfile[11][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y35_N19
dffeas \rfile[9][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][1] .is_wysiwyg = "true";
defparam \rfile[9][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N9
dffeas \rfile[10][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][1] .is_wysiwyg = "true";
defparam \rfile[10][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N15
dffeas \rfile[8][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][1] .is_wysiwyg = "true";
defparam \rfile[8][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N14
cycloneive_lcell_comb \Mux30~10 (
// Equation(s):
// \Mux30~10_combout  = (instruction_D[22] & ((\rfile[10][1]~q ) # ((instruction_D[21])))) # (!instruction_D[22] & (((\rfile[8][1]~q  & !instruction_D[21]))))

	.dataa(instruction_D_22),
	.datab(\rfile[10][1]~q ),
	.datac(\rfile[8][1]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux30~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~10 .lut_mask = 16'hAAD8;
defparam \Mux30~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N18
cycloneive_lcell_comb \Mux30~11 (
// Equation(s):
// \Mux30~11_combout  = (instruction_D[21] & ((\Mux30~10_combout  & (\rfile[11][1]~q )) # (!\Mux30~10_combout  & ((\rfile[9][1]~q ))))) # (!instruction_D[21] & (((\Mux30~10_combout ))))

	.dataa(\rfile[11][1]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[9][1]~q ),
	.datad(\Mux30~10_combout ),
	.cin(gnd),
	.combout(\Mux30~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~11 .lut_mask = 16'hBBC0;
defparam \Mux30~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N9
dffeas \rfile[15][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][1] .is_wysiwyg = "true";
defparam \rfile[15][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y33_N25
dffeas \rfile[14][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][1] .is_wysiwyg = "true";
defparam \rfile[14][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N6
cycloneive_lcell_comb \rfile[13][1]~feeder (
// Equation(s):
// \rfile[13][1]~feeder_combout  = \wdat_WB[1]~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[13][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[13][1]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[13][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N7
dffeas \rfile[13][1] (
	.clk(!CLK),
	.d(\rfile[13][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][1] .is_wysiwyg = "true";
defparam \rfile[13][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N28
cycloneive_lcell_comb \Mux30~17 (
// Equation(s):
// \Mux30~17_combout  = (instruction_D[21] & (((instruction_D[22]) # (\rfile[13][1]~q )))) # (!instruction_D[21] & (\rfile[12][1]~q  & (!instruction_D[22])))

	.dataa(\rfile[12][1]~q ),
	.datab(instruction_D_21),
	.datac(instruction_D_22),
	.datad(\rfile[13][1]~q ),
	.cin(gnd),
	.combout(\Mux30~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~17 .lut_mask = 16'hCEC2;
defparam \Mux30~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N18
cycloneive_lcell_comb \Mux30~18 (
// Equation(s):
// \Mux30~18_combout  = (instruction_D[22] & ((\Mux30~17_combout  & (\rfile[15][1]~q )) # (!\Mux30~17_combout  & ((\rfile[14][1]~q ))))) # (!instruction_D[22] & (((\Mux30~17_combout ))))

	.dataa(\rfile[15][1]~q ),
	.datab(\rfile[14][1]~q ),
	.datac(instruction_D_22),
	.datad(\Mux30~17_combout ),
	.cin(gnd),
	.combout(\Mux30~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~18 .lut_mask = 16'hAFC0;
defparam \Mux30~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N8
cycloneive_lcell_comb \rfile[7][1]~feeder (
// Equation(s):
// \rfile[7][1]~feeder_combout  = \wdat_WB[1]~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_1),
	.cin(gnd),
	.combout(\rfile[7][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[7][1]~feeder .lut_mask = 16'hFF00;
defparam \rfile[7][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N9
dffeas \rfile[7][1] (
	.clk(!CLK),
	.d(\rfile[7][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][1] .is_wysiwyg = "true";
defparam \rfile[7][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y36_N5
dffeas \rfile[6][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][1] .is_wysiwyg = "true";
defparam \rfile[6][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N4
cycloneive_lcell_comb \Mux30~13 (
// Equation(s):
// \Mux30~13_combout  = (\Mux30~12_combout  & ((\rfile[7][1]~q ) # ((!instruction_D[22])))) # (!\Mux30~12_combout  & (((\rfile[6][1]~q  & instruction_D[22]))))

	.dataa(\Mux30~12_combout ),
	.datab(\rfile[7][1]~q ),
	.datac(\rfile[6][1]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux30~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~13 .lut_mask = 16'hD8AA;
defparam \Mux30~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y34_N19
dffeas \rfile[1][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][1] .is_wysiwyg = "true";
defparam \rfile[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y34_N29
dffeas \rfile[3][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][1] .is_wysiwyg = "true";
defparam \rfile[3][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N18
cycloneive_lcell_comb \Mux30~14 (
// Equation(s):
// \Mux30~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][1]~q ))) # (!instruction_D[22] & (\rfile[1][1]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][1]~q ),
	.datad(\rfile[3][1]~q ),
	.cin(gnd),
	.combout(\Mux30~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~14 .lut_mask = 16'hC840;
defparam \Mux30~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N20
cycloneive_lcell_comb \Mux30~15 (
// Equation(s):
// \Mux30~15_combout  = (\Mux30~14_combout ) # ((\rfile[2][1]~q  & (!instruction_D[21] & instruction_D[22])))

	.dataa(\rfile[2][1]~q ),
	.datab(instruction_D_21),
	.datac(instruction_D_22),
	.datad(\Mux30~14_combout ),
	.cin(gnd),
	.combout(\Mux30~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~15 .lut_mask = 16'hFF20;
defparam \Mux30~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N18
cycloneive_lcell_comb \Mux30~16 (
// Equation(s):
// \Mux30~16_combout  = (instruction_D[24] & (((instruction_D[23])))) # (!instruction_D[24] & ((instruction_D[23] & (\Mux30~13_combout )) # (!instruction_D[23] & ((\Mux30~15_combout )))))

	.dataa(instruction_D_24),
	.datab(\Mux30~13_combout ),
	.datac(instruction_D_23),
	.datad(\Mux30~15_combout ),
	.cin(gnd),
	.combout(\Mux30~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~16 .lut_mask = 16'hE5E0;
defparam \Mux30~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N11
dffeas \rfile[29][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][0] .is_wysiwyg = "true";
defparam \rfile[29][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N17
dffeas \rfile[21][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][0] .is_wysiwyg = "true";
defparam \rfile[21][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N21
dffeas \rfile[25][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][0] .is_wysiwyg = "true";
defparam \rfile[25][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N3
dffeas \rfile[17][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][0] .is_wysiwyg = "true";
defparam \rfile[17][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N20
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[25][0]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[17][0]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[25][0]~q ),
	.datad(\rfile[17][0]~q ),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'hB9A8;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N16
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (instruction_D[18] & ((\Mux63~0_combout  & (\rfile[29][0]~q )) # (!\Mux63~0_combout  & ((\rfile[21][0]~q ))))) # (!instruction_D[18] & (((\Mux63~0_combout ))))

	.dataa(\rfile[29][0]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[21][0]~q ),
	.datad(\Mux63~0_combout ),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'hBBC0;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y31_N9
dffeas \rfile[23][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][0] .is_wysiwyg = "true";
defparam \rfile[23][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y31_N11
dffeas \rfile[31][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][0] .is_wysiwyg = "true";
defparam \rfile[31][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N25
dffeas \rfile[27][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][0] .is_wysiwyg = "true";
defparam \rfile[27][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N7
dffeas \rfile[19][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][0] .is_wysiwyg = "true";
defparam \rfile[19][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N24
cycloneive_lcell_comb \Mux63~7 (
// Equation(s):
// \Mux63~7_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[27][0]~q )) # (!instruction_D[19] & ((\rfile[19][0]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[27][0]~q ),
	.datad(\rfile[19][0]~q ),
	.cin(gnd),
	.combout(\Mux63~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~7 .lut_mask = 16'hD9C8;
defparam \Mux63~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N10
cycloneive_lcell_comb \Mux63~8 (
// Equation(s):
// \Mux63~8_combout  = (instruction_D[18] & ((\Mux63~7_combout  & ((\rfile[31][0]~q ))) # (!\Mux63~7_combout  & (\rfile[23][0]~q )))) # (!instruction_D[18] & (((\Mux63~7_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[23][0]~q ),
	.datac(\rfile[31][0]~q ),
	.datad(\Mux63~7_combout ),
	.cin(gnd),
	.combout(\Mux63~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~8 .lut_mask = 16'hF588;
defparam \Mux63~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y34_N13
dffeas \rfile[18][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][0] .is_wysiwyg = "true";
defparam \rfile[18][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y34_N3
dffeas \rfile[22][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][0] .is_wysiwyg = "true";
defparam \rfile[22][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N12
cycloneive_lcell_comb \Mux63~2 (
// Equation(s):
// \Mux63~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[22][0]~q ))) # (!instruction_D[18] & (\rfile[18][0]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][0]~q ),
	.datad(\rfile[22][0]~q ),
	.cin(gnd),
	.combout(\Mux63~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~2 .lut_mask = 16'hDC98;
defparam \Mux63~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y34_N9
dffeas \rfile[30][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][0] .is_wysiwyg = "true";
defparam \rfile[30][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y34_N7
dffeas \rfile[26][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][0] .is_wysiwyg = "true";
defparam \rfile[26][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N8
cycloneive_lcell_comb \Mux63~3 (
// Equation(s):
// \Mux63~3_combout  = (instruction_D[19] & ((\Mux63~2_combout  & (\rfile[30][0]~q )) # (!\Mux63~2_combout  & ((\rfile[26][0]~q ))))) # (!instruction_D[19] & (\Mux63~2_combout ))

	.dataa(instruction_D_19),
	.datab(\Mux63~2_combout ),
	.datac(\rfile[30][0]~q ),
	.datad(\rfile[26][0]~q ),
	.cin(gnd),
	.combout(\Mux63~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~3 .lut_mask = 16'hE6C4;
defparam \Mux63~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N13
dffeas \rfile[24][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][0] .is_wysiwyg = "true";
defparam \rfile[24][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y31_N23
dffeas \rfile[20][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][0] .is_wysiwyg = "true";
defparam \rfile[20][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y31_N1
dffeas \rfile[16][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][0] .is_wysiwyg = "true";
defparam \rfile[16][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N22
cycloneive_lcell_comb \Mux63~4 (
// Equation(s):
// \Mux63~4_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[20][0]~q )))) # (!instruction_D[18] & (!instruction_D[19] & ((\rfile[16][0]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[20][0]~q ),
	.datad(\rfile[16][0]~q ),
	.cin(gnd),
	.combout(\Mux63~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~4 .lut_mask = 16'hB9A8;
defparam \Mux63~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N12
cycloneive_lcell_comb \Mux63~5 (
// Equation(s):
// \Mux63~5_combout  = (instruction_D[19] & ((\Mux63~4_combout  & (\rfile[28][0]~q )) # (!\Mux63~4_combout  & ((\rfile[24][0]~q ))))) # (!instruction_D[19] & (((\Mux63~4_combout ))))

	.dataa(\rfile[28][0]~q ),
	.datab(instruction_D_19),
	.datac(\rfile[24][0]~q ),
	.datad(\Mux63~4_combout ),
	.cin(gnd),
	.combout(\Mux63~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~5 .lut_mask = 16'hBBC0;
defparam \Mux63~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N0
cycloneive_lcell_comb \Mux63~6 (
// Equation(s):
// \Mux63~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\Mux63~3_combout )) # (!instruction_D[17] & ((\Mux63~5_combout )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux63~3_combout ),
	.datad(\Mux63~5_combout ),
	.cin(gnd),
	.combout(\Mux63~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~6 .lut_mask = 16'hD9C8;
defparam \Mux63~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N21
dffeas \rfile[3][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][0] .is_wysiwyg = "true";
defparam \rfile[3][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N19
dffeas \rfile[1][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][0] .is_wysiwyg = "true";
defparam \rfile[1][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N20
cycloneive_lcell_comb \Mux63~14 (
// Equation(s):
// \Mux63~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][0]~q )) # (!instruction_D[17] & ((\rfile[1][0]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[3][0]~q ),
	.datad(\rfile[1][0]~q ),
	.cin(gnd),
	.combout(\Mux63~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~14 .lut_mask = 16'hC480;
defparam \Mux63~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N16
cycloneive_lcell_comb \rfile[2][0]~feeder (
// Equation(s):
// \rfile[2][0]~feeder_combout  = \wdat_WB[0]~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_0),
	.cin(gnd),
	.combout(\rfile[2][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][0]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N17
dffeas \rfile[2][0] (
	.clk(!CLK),
	.d(\rfile[2][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][0] .is_wysiwyg = "true";
defparam \rfile[2][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N26
cycloneive_lcell_comb \Mux63~15 (
// Equation(s):
// \Mux63~15_combout  = (\Mux63~14_combout ) # ((!instruction_D[16] & (instruction_D[17] & \rfile[2][0]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux63~14_combout ),
	.datad(\rfile[2][0]~q ),
	.cin(gnd),
	.combout(\Mux63~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~15 .lut_mask = 16'hF4F0;
defparam \Mux63~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N5
dffeas \rfile[11][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][0] .is_wysiwyg = "true";
defparam \rfile[11][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y35_N7
dffeas \rfile[9][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][0] .is_wysiwyg = "true";
defparam \rfile[9][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N1
dffeas \rfile[10][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][0] .is_wysiwyg = "true";
defparam \rfile[10][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N15
dffeas \rfile[8][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][0] .is_wysiwyg = "true";
defparam \rfile[8][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N0
cycloneive_lcell_comb \Mux63~12 (
// Equation(s):
// \Mux63~12_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\rfile[10][0]~q )))) # (!instruction_D[17] & (!instruction_D[16] & ((\rfile[8][0]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[10][0]~q ),
	.datad(\rfile[8][0]~q ),
	.cin(gnd),
	.combout(\Mux63~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~12 .lut_mask = 16'hB9A8;
defparam \Mux63~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N6
cycloneive_lcell_comb \Mux63~13 (
// Equation(s):
// \Mux63~13_combout  = (instruction_D[16] & ((\Mux63~12_combout  & (\rfile[11][0]~q )) # (!\Mux63~12_combout  & ((\rfile[9][0]~q ))))) # (!instruction_D[16] & (((\Mux63~12_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][0]~q ),
	.datac(\rfile[9][0]~q ),
	.datad(\Mux63~12_combout ),
	.cin(gnd),
	.combout(\Mux63~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~13 .lut_mask = 16'hDDA0;
defparam \Mux63~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N12
cycloneive_lcell_comb \Mux63~16 (
// Equation(s):
// \Mux63~16_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\Mux63~13_combout )))) # (!instruction_D[19] & (!instruction_D[18] & (\Mux63~15_combout )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux63~15_combout ),
	.datad(\Mux63~13_combout ),
	.cin(gnd),
	.combout(\Mux63~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~16 .lut_mask = 16'hBA98;
defparam \Mux63~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N29
dffeas \rfile[13][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][0] .is_wysiwyg = "true";
defparam \rfile[13][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N28
cycloneive_lcell_comb \Mux63~17 (
// Equation(s):
// \Mux63~17_combout  = (instruction_D[16] & (((\rfile[13][0]~q ) # (instruction_D[17])))) # (!instruction_D[16] & (\rfile[12][0]~q  & ((!instruction_D[17]))))

	.dataa(\rfile[12][0]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[13][0]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux63~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~17 .lut_mask = 16'hCCE2;
defparam \Mux63~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N1
dffeas \rfile[14][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][0] .is_wysiwyg = "true";
defparam \rfile[14][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N27
dffeas \rfile[15][0] (
	.clk(!CLK),
	.d(wdat_WB_0),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][0] .is_wysiwyg = "true";
defparam \rfile[15][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N0
cycloneive_lcell_comb \Mux63~18 (
// Equation(s):
// \Mux63~18_combout  = (instruction_D[17] & ((\Mux63~17_combout  & ((\rfile[15][0]~q ))) # (!\Mux63~17_combout  & (\rfile[14][0]~q )))) # (!instruction_D[17] & (\Mux63~17_combout ))

	.dataa(instruction_D_17),
	.datab(\Mux63~17_combout ),
	.datac(\rfile[14][0]~q ),
	.datad(\rfile[15][0]~q ),
	.cin(gnd),
	.combout(\Mux63~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~18 .lut_mask = 16'hEC64;
defparam \Mux63~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N31
dffeas \rfile[7][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][0] .is_wysiwyg = "true";
defparam \rfile[7][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N1
dffeas \rfile[6][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][0] .is_wysiwyg = "true";
defparam \rfile[6][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N19
dffeas \rfile[5][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][0] .is_wysiwyg = "true";
defparam \rfile[5][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y28_N15
dffeas \rfile[4][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][0] .is_wysiwyg = "true";
defparam \rfile[4][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N18
cycloneive_lcell_comb \Mux63~10 (
// Equation(s):
// \Mux63~10_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[5][0]~q )) # (!instruction_D[16] & ((\rfile[4][0]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[5][0]~q ),
	.datad(\rfile[4][0]~q ),
	.cin(gnd),
	.combout(\Mux63~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~10 .lut_mask = 16'hD9C8;
defparam \Mux63~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N0
cycloneive_lcell_comb \Mux63~11 (
// Equation(s):
// \Mux63~11_combout  = (instruction_D[17] & ((\Mux63~10_combout  & (\rfile[7][0]~q )) # (!\Mux63~10_combout  & ((\rfile[6][0]~q ))))) # (!instruction_D[17] & (((\Mux63~10_combout ))))

	.dataa(\rfile[7][0]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[6][0]~q ),
	.datad(\Mux63~10_combout ),
	.cin(gnd),
	.combout(\Mux63~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~11 .lut_mask = 16'hBBC0;
defparam \Mux63~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N27
dffeas \rfile[21][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][1] .is_wysiwyg = "true";
defparam \rfile[21][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N26
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[21][1]~q )))) # (!instruction_D[18] & (!instruction_D[19] & ((\rfile[17][1]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[21][1]~q ),
	.datad(\rfile[17][1]~q ),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'hB9A8;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N0
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (instruction_D[19] & ((\Mux62~0_combout  & (\rfile[29][1]~q )) # (!\Mux62~0_combout  & ((\rfile[25][1]~q ))))) # (!instruction_D[19] & (((\Mux62~0_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[29][1]~q ),
	.datac(\rfile[25][1]~q ),
	.datad(\Mux62~0_combout ),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'hDDA0;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N26
cycloneive_lcell_comb \Mux62~4 (
// Equation(s):
// \Mux62~4_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[24][1]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[16][1]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[24][1]~q ),
	.datad(\rfile[16][1]~q ),
	.cin(gnd),
	.combout(\Mux62~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~4 .lut_mask = 16'hB9A8;
defparam \Mux62~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N10
cycloneive_lcell_comb \Mux62~5 (
// Equation(s):
// \Mux62~5_combout  = (instruction_D[18] & ((\Mux62~4_combout  & ((\rfile[28][1]~q ))) # (!\Mux62~4_combout  & (\rfile[20][1]~q )))) # (!instruction_D[18] & (((\Mux62~4_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[20][1]~q ),
	.datac(\Mux62~4_combout ),
	.datad(\rfile[28][1]~q ),
	.cin(gnd),
	.combout(\Mux62~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~5 .lut_mask = 16'hF858;
defparam \Mux62~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N24
cycloneive_lcell_comb \Mux62~3 (
// Equation(s):
// \Mux62~3_combout  = (\Mux62~2_combout  & (((\rfile[30][1]~q ) # (!instruction_D[18])))) # (!\Mux62~2_combout  & (\rfile[22][1]~q  & ((instruction_D[18]))))

	.dataa(\Mux62~2_combout ),
	.datab(\rfile[22][1]~q ),
	.datac(\rfile[30][1]~q ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux62~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~3 .lut_mask = 16'hE4AA;
defparam \Mux62~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N4
cycloneive_lcell_comb \Mux62~6 (
// Equation(s):
// \Mux62~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\Mux62~3_combout ))) # (!instruction_D[17] & (\Mux62~5_combout ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux62~5_combout ),
	.datad(\Mux62~3_combout ),
	.cin(gnd),
	.combout(\Mux62~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~6 .lut_mask = 16'hDC98;
defparam \Mux62~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N0
cycloneive_lcell_comb \Mux62~7 (
// Equation(s):
// \Mux62~7_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[23][1]~q )) # (!instruction_D[18] & ((\rfile[19][1]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[23][1]~q ),
	.datad(\rfile[19][1]~q ),
	.cin(gnd),
	.combout(\Mux62~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~7 .lut_mask = 16'hD9C8;
defparam \Mux62~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N8
cycloneive_lcell_comb \Mux62~8 (
// Equation(s):
// \Mux62~8_combout  = (instruction_D[19] & ((\Mux62~7_combout  & (\rfile[31][1]~q )) # (!\Mux62~7_combout  & ((\rfile[27][1]~q ))))) # (!instruction_D[19] & (((\Mux62~7_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[31][1]~q ),
	.datac(\rfile[27][1]~q ),
	.datad(\Mux62~7_combout ),
	.cin(gnd),
	.combout(\Mux62~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~8 .lut_mask = 16'hDDA0;
defparam \Mux62~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N8
cycloneive_lcell_comb \Mux62~10 (
// Equation(s):
// \Mux62~10_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][1]~q ))) # (!instruction_D[17] & (\rfile[8][1]~q ))))

	.dataa(instruction_D_16),
	.datab(\rfile[8][1]~q ),
	.datac(\rfile[10][1]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux62~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~10 .lut_mask = 16'hFA44;
defparam \Mux62~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N12
cycloneive_lcell_comb \Mux62~11 (
// Equation(s):
// \Mux62~11_combout  = (instruction_D[16] & ((\Mux62~10_combout  & ((\rfile[11][1]~q ))) # (!\Mux62~10_combout  & (\rfile[9][1]~q )))) # (!instruction_D[16] & (((\Mux62~10_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[9][1]~q ),
	.datac(\rfile[11][1]~q ),
	.datad(\Mux62~10_combout ),
	.cin(gnd),
	.combout(\Mux62~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~11 .lut_mask = 16'hF588;
defparam \Mux62~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N10
cycloneive_lcell_comb \Mux62~17 (
// Equation(s):
// \Mux62~17_combout  = (instruction_D[17] & (((instruction_D[16])))) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[13][1]~q ))) # (!instruction_D[16] & (\rfile[12][1]~q ))))

	.dataa(\rfile[12][1]~q ),
	.datab(instruction_D_17),
	.datac(instruction_D_16),
	.datad(\rfile[13][1]~q ),
	.cin(gnd),
	.combout(\Mux62~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~17 .lut_mask = 16'hF2C2;
defparam \Mux62~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N24
cycloneive_lcell_comb \Mux62~18 (
// Equation(s):
// \Mux62~18_combout  = (instruction_D[17] & ((\Mux62~17_combout  & (\rfile[15][1]~q )) # (!\Mux62~17_combout  & ((\rfile[14][1]~q ))))) # (!instruction_D[17] & (((\Mux62~17_combout ))))

	.dataa(\rfile[15][1]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[14][1]~q ),
	.datad(\Mux62~17_combout ),
	.cin(gnd),
	.combout(\Mux62~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~18 .lut_mask = 16'hBBC0;
defparam \Mux62~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N28
cycloneive_lcell_comb \Mux62~14 (
// Equation(s):
// \Mux62~14_combout  = (instruction_D[16] & ((instruction_D[17] & (\rfile[3][1]~q )) # (!instruction_D[17] & ((\rfile[1][1]~q )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[3][1]~q ),
	.datad(\rfile[1][1]~q ),
	.cin(gnd),
	.combout(\Mux62~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~14 .lut_mask = 16'hA280;
defparam \Mux62~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N30
cycloneive_lcell_comb \Mux62~15 (
// Equation(s):
// \Mux62~15_combout  = (\Mux62~14_combout ) # ((\rfile[2][1]~q  & (instruction_D[17] & !instruction_D[16])))

	.dataa(\rfile[2][1]~q ),
	.datab(instruction_D_17),
	.datac(instruction_D_16),
	.datad(\Mux62~14_combout ),
	.cin(gnd),
	.combout(\Mux62~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~15 .lut_mask = 16'hFF08;
defparam \Mux62~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N9
dffeas \rfile[5][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][1] .is_wysiwyg = "true";
defparam \rfile[5][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N8
cycloneive_lcell_comb \Mux62~12 (
// Equation(s):
// \Mux62~12_combout  = (instruction_D[16] & (((\rfile[5][1]~q ) # (instruction_D[17])))) # (!instruction_D[16] & (\rfile[4][1]~q  & ((!instruction_D[17]))))

	.dataa(\rfile[4][1]~q ),
	.datab(instruction_D_16),
	.datac(\rfile[5][1]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux62~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~12 .lut_mask = 16'hCCE2;
defparam \Mux62~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N24
cycloneive_lcell_comb \Mux62~13 (
// Equation(s):
// \Mux62~13_combout  = (instruction_D[17] & ((\Mux62~12_combout  & (\rfile[7][1]~q )) # (!\Mux62~12_combout  & ((\rfile[6][1]~q ))))) # (!instruction_D[17] & (((\Mux62~12_combout ))))

	.dataa(\rfile[7][1]~q ),
	.datab(\rfile[6][1]~q ),
	.datac(instruction_D_17),
	.datad(\Mux62~12_combout ),
	.cin(gnd),
	.combout(\Mux62~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~13 .lut_mask = 16'hAFC0;
defparam \Mux62~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N28
cycloneive_lcell_comb \Mux62~16 (
// Equation(s):
// \Mux62~16_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\Mux62~13_combout ))) # (!instruction_D[18] & (\Mux62~15_combout ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux62~15_combout ),
	.datad(\Mux62~13_combout ),
	.cin(gnd),
	.combout(\Mux62~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~16 .lut_mask = 16'hDC98;
defparam \Mux62~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N3
dffeas \rfile[23][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][4] .is_wysiwyg = "true";
defparam \rfile[23][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N21
dffeas \rfile[31][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][4] .is_wysiwyg = "true";
defparam \rfile[31][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N21
dffeas \rfile[27][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][4] .is_wysiwyg = "true";
defparam \rfile[27][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N3
dffeas \rfile[19][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][4] .is_wysiwyg = "true";
defparam \rfile[19][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N20
cycloneive_lcell_comb \Mux27~7 (
// Equation(s):
// \Mux27~7_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[27][4]~q )) # (!instruction_D[24] & ((\rfile[19][4]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[27][4]~q ),
	.datad(\rfile[19][4]~q ),
	.cin(gnd),
	.combout(\Mux27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~7 .lut_mask = 16'hD9C8;
defparam \Mux27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N20
cycloneive_lcell_comb \Mux27~8 (
// Equation(s):
// \Mux27~8_combout  = (instruction_D[23] & ((\Mux27~7_combout  & ((\rfile[31][4]~q ))) # (!\Mux27~7_combout  & (\rfile[23][4]~q )))) # (!instruction_D[23] & (((\Mux27~7_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[23][4]~q ),
	.datac(\rfile[31][4]~q ),
	.datad(\Mux27~7_combout ),
	.cin(gnd),
	.combout(\Mux27~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~8 .lut_mask = 16'hF588;
defparam \Mux27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N9
dffeas \rfile[25][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][4] .is_wysiwyg = "true";
defparam \rfile[25][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N6
cycloneive_lcell_comb \rfile[17][4]~feeder (
// Equation(s):
// \rfile[17][4]~feeder_combout  = \wdat_WB[4]~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[17][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[17][4]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[17][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N7
dffeas \rfile[17][4] (
	.clk(!CLK),
	.d(\rfile[17][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][4] .is_wysiwyg = "true";
defparam \rfile[17][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N30
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[25][4]~q )) # (!instruction_D[24] & ((\rfile[17][4]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[25][4]~q ),
	.datad(\rfile[17][4]~q ),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hD9C8;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N7
dffeas \rfile[21][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][4] .is_wysiwyg = "true";
defparam \rfile[21][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N13
dffeas \rfile[29][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][4] .is_wysiwyg = "true";
defparam \rfile[29][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N6
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (\Mux27~0_combout  & (((\rfile[29][4]~q )) # (!instruction_D[23]))) # (!\Mux27~0_combout  & (instruction_D[23] & (\rfile[21][4]~q )))

	.dataa(\Mux27~0_combout ),
	.datab(instruction_D_23),
	.datac(\rfile[21][4]~q ),
	.datad(\rfile[29][4]~q ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hEA62;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y34_N4
cycloneive_lcell_comb \rfile[26][4]~feeder (
// Equation(s):
// \rfile[26][4]~feeder_combout  = \wdat_WB[4]~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_4),
	.cin(gnd),
	.combout(\rfile[26][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[26][4]~feeder .lut_mask = 16'hFF00;
defparam \rfile[26][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y34_N5
dffeas \rfile[26][4] (
	.clk(!CLK),
	.d(\rfile[26][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][4] .is_wysiwyg = "true";
defparam \rfile[26][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N14
cycloneive_lcell_comb \rfile[22][4]~feeder (
// Equation(s):
// \rfile[22][4]~feeder_combout  = \wdat_WB[4]~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[22][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[22][4]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[22][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y34_N15
dffeas \rfile[22][4] (
	.clk(!CLK),
	.d(\rfile[22][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][4] .is_wysiwyg = "true";
defparam \rfile[22][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y34_N21
dffeas \rfile[18][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][4] .is_wysiwyg = "true";
defparam \rfile[18][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N10
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[22][4]~q )) # (!instruction_D[23] & ((\rfile[18][4]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[22][4]~q ),
	.datad(\rfile[18][4]~q ),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'hD9C8;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y34_N24
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (instruction_D[24] & ((\Mux27~2_combout  & (\rfile[30][4]~q )) # (!\Mux27~2_combout  & ((\rfile[26][4]~q ))))) # (!instruction_D[24] & (((\Mux27~2_combout ))))

	.dataa(\rfile[30][4]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[26][4]~q ),
	.datad(\Mux27~2_combout ),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'hBBC0;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N17
dffeas \rfile[24][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][4] .is_wysiwyg = "true";
defparam \rfile[24][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N3
dffeas \rfile[28][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][4] .is_wysiwyg = "true";
defparam \rfile[28][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y32_N5
dffeas \rfile[20][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][4] .is_wysiwyg = "true";
defparam \rfile[20][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N10
cycloneive_lcell_comb \rfile[16][4]~feeder (
// Equation(s):
// \rfile[16][4]~feeder_combout  = \wdat_WB[4]~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[16][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[16][4]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[16][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y32_N11
dffeas \rfile[16][4] (
	.clk(!CLK),
	.d(\rfile[16][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][4] .is_wysiwyg = "true";
defparam \rfile[16][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N0
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[20][4]~q )) # (!instruction_D[23] & ((\rfile[16][4]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[20][4]~q ),
	.datad(\rfile[16][4]~q ),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'hD9C8;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N2
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// \Mux27~5_combout  = (instruction_D[24] & ((\Mux27~4_combout  & ((\rfile[28][4]~q ))) # (!\Mux27~4_combout  & (\rfile[24][4]~q )))) # (!instruction_D[24] & (((\Mux27~4_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[24][4]~q ),
	.datac(\rfile[28][4]~q ),
	.datad(\Mux27~4_combout ),
	.cin(gnd),
	.combout(\Mux27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hF588;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N2
cycloneive_lcell_comb \Mux27~6 (
// Equation(s):
// \Mux27~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\Mux27~3_combout )) # (!instruction_D[22] & ((\Mux27~5_combout )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux27~3_combout ),
	.datad(\Mux27~5_combout ),
	.cin(gnd),
	.combout(\Mux27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~6 .lut_mask = 16'hD9C8;
defparam \Mux27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N23
dffeas \rfile[15][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][4] .is_wysiwyg = "true";
defparam \rfile[15][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N7
dffeas \rfile[14][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][4] .is_wysiwyg = "true";
defparam \rfile[14][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N1
dffeas \rfile[13][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][4] .is_wysiwyg = "true";
defparam \rfile[13][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N3
dffeas \rfile[12][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][4] .is_wysiwyg = "true";
defparam \rfile[12][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N0
cycloneive_lcell_comb \Mux27~17 (
// Equation(s):
// \Mux27~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][4]~q )) # (!instruction_D[21] & ((\rfile[12][4]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[13][4]~q ),
	.datad(\rfile[12][4]~q ),
	.cin(gnd),
	.combout(\Mux27~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~17 .lut_mask = 16'hD9C8;
defparam \Mux27~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N6
cycloneive_lcell_comb \Mux27~18 (
// Equation(s):
// \Mux27~18_combout  = (instruction_D[22] & ((\Mux27~17_combout  & (\rfile[15][4]~q )) # (!\Mux27~17_combout  & ((\rfile[14][4]~q ))))) # (!instruction_D[22] & (((\Mux27~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[15][4]~q ),
	.datac(\rfile[14][4]~q ),
	.datad(\Mux27~17_combout ),
	.cin(gnd),
	.combout(\Mux27~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~18 .lut_mask = 16'hDDA0;
defparam \Mux27~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N15
dffeas \rfile[7][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][4] .is_wysiwyg = "true";
defparam \rfile[7][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N25
dffeas \rfile[6][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][4] .is_wysiwyg = "true";
defparam \rfile[6][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N17
dffeas \rfile[5][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][4] .is_wysiwyg = "true";
defparam \rfile[5][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N7
dffeas \rfile[4][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][4] .is_wysiwyg = "true";
defparam \rfile[4][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N16
cycloneive_lcell_comb \Mux27~10 (
// Equation(s):
// \Mux27~10_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[5][4]~q )) # (!instruction_D[21] & ((\rfile[4][4]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[5][4]~q ),
	.datad(\rfile[4][4]~q ),
	.cin(gnd),
	.combout(\Mux27~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~10 .lut_mask = 16'hD9C8;
defparam \Mux27~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N24
cycloneive_lcell_comb \Mux27~11 (
// Equation(s):
// \Mux27~11_combout  = (instruction_D[22] & ((\Mux27~10_combout  & (\rfile[7][4]~q )) # (!\Mux27~10_combout  & ((\rfile[6][4]~q ))))) # (!instruction_D[22] & (((\Mux27~10_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[7][4]~q ),
	.datac(\rfile[6][4]~q ),
	.datad(\Mux27~10_combout ),
	.cin(gnd),
	.combout(\Mux27~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~11 .lut_mask = 16'hDDA0;
defparam \Mux27~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N3
dffeas \rfile[3][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][4] .is_wysiwyg = "true";
defparam \rfile[3][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N29
dffeas \rfile[1][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][4] .is_wysiwyg = "true";
defparam \rfile[1][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N2
cycloneive_lcell_comb \Mux27~14 (
// Equation(s):
// \Mux27~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][4]~q )) # (!instruction_D[22] & ((\rfile[1][4]~q )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[3][4]~q ),
	.datad(\rfile[1][4]~q ),
	.cin(gnd),
	.combout(\Mux27~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~14 .lut_mask = 16'hA280;
defparam \Mux27~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N8
cycloneive_lcell_comb \rfile[2][4]~feeder (
// Equation(s):
// \rfile[2][4]~feeder_combout  = \wdat_WB[4]~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_4),
	.cin(gnd),
	.combout(\rfile[2][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][4]~feeder .lut_mask = 16'hFF00;
defparam \rfile[2][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N9
dffeas \rfile[2][4] (
	.clk(!CLK),
	.d(\rfile[2][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][4] .is_wysiwyg = "true";
defparam \rfile[2][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N30
cycloneive_lcell_comb \Mux27~15 (
// Equation(s):
// \Mux27~15_combout  = (\Mux27~14_combout ) # ((!instruction_D[21] & (instruction_D[22] & \rfile[2][4]~q )))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux27~14_combout ),
	.datad(\rfile[2][4]~q ),
	.cin(gnd),
	.combout(\Mux27~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~15 .lut_mask = 16'hF4F0;
defparam \Mux27~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N2
cycloneive_lcell_comb \rfile[11][4]~feeder (
// Equation(s):
// \rfile[11][4]~feeder_combout  = \wdat_WB[4]~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_4),
	.cin(gnd),
	.combout(\rfile[11][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][4]~feeder .lut_mask = 16'hFF00;
defparam \rfile[11][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N3
dffeas \rfile[11][4] (
	.clk(!CLK),
	.d(\rfile[11][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][4] .is_wysiwyg = "true";
defparam \rfile[11][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N29
dffeas \rfile[9][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][4] .is_wysiwyg = "true";
defparam \rfile[9][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N25
dffeas \rfile[10][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][4] .is_wysiwyg = "true";
defparam \rfile[10][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N3
dffeas \rfile[8][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][4] .is_wysiwyg = "true";
defparam \rfile[8][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N24
cycloneive_lcell_comb \Mux27~12 (
// Equation(s):
// \Mux27~12_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][4]~q )))) # (!instruction_D[22] & (!instruction_D[21] & ((\rfile[8][4]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[10][4]~q ),
	.datad(\rfile[8][4]~q ),
	.cin(gnd),
	.combout(\Mux27~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~12 .lut_mask = 16'hB9A8;
defparam \Mux27~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N28
cycloneive_lcell_comb \Mux27~13 (
// Equation(s):
// \Mux27~13_combout  = (instruction_D[21] & ((\Mux27~12_combout  & (\rfile[11][4]~q )) # (!\Mux27~12_combout  & ((\rfile[9][4]~q ))))) # (!instruction_D[21] & (((\Mux27~12_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[11][4]~q ),
	.datac(\rfile[9][4]~q ),
	.datad(\Mux27~12_combout ),
	.cin(gnd),
	.combout(\Mux27~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~13 .lut_mask = 16'hDDA0;
defparam \Mux27~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N28
cycloneive_lcell_comb \Mux27~16 (
// Equation(s):
// \Mux27~16_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\Mux27~13_combout ))) # (!instruction_D[24] & (\Mux27~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux27~15_combout ),
	.datad(\Mux27~13_combout ),
	.cin(gnd),
	.combout(\Mux27~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~16 .lut_mask = 16'hDC98;
defparam \Mux27~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N20
cycloneive_lcell_comb \rfile[23][3]~feeder (
// Equation(s):
// \rfile[23][3]~feeder_combout  = \wdat_WB[3]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[23][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[23][3]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[23][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y29_N21
dffeas \rfile[23][3] (
	.clk(!CLK),
	.d(\rfile[23][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[23][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[23][3] .is_wysiwyg = "true";
defparam \rfile[23][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y29_N11
dffeas \rfile[31][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[31][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[31][3] .is_wysiwyg = "true";
defparam \rfile[31][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y29_N9
dffeas \rfile[27][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[27][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[27][3] .is_wysiwyg = "true";
defparam \rfile[27][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N8
cycloneive_lcell_comb \Mux28~7 (
// Equation(s):
// \Mux28~7_combout  = (instruction_D[24] & (((\rfile[27][3]~q ) # (instruction_D[23])))) # (!instruction_D[24] & (\rfile[19][3]~q  & ((!instruction_D[23]))))

	.dataa(\rfile[19][3]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[27][3]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~7 .lut_mask = 16'hCCE2;
defparam \Mux28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N10
cycloneive_lcell_comb \Mux28~8 (
// Equation(s):
// \Mux28~8_combout  = (instruction_D[23] & ((\Mux28~7_combout  & ((\rfile[31][3]~q ))) # (!\Mux28~7_combout  & (\rfile[23][3]~q )))) # (!instruction_D[23] & (((\Mux28~7_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[23][3]~q ),
	.datac(\rfile[31][3]~q ),
	.datad(\Mux28~7_combout ),
	.cin(gnd),
	.combout(\Mux28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~8 .lut_mask = 16'hF588;
defparam \Mux28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N26
cycloneive_lcell_comb \rfile[21][3]~feeder (
// Equation(s):
// \rfile[21][3]~feeder_combout  = \wdat_WB[3]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_3),
	.cin(gnd),
	.combout(\rfile[21][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[21][3]~feeder .lut_mask = 16'hFF00;
defparam \rfile[21][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N27
dffeas \rfile[21][3] (
	.clk(!CLK),
	.d(\rfile[21][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[21][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[21][3] .is_wysiwyg = "true";
defparam \rfile[21][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N24
cycloneive_lcell_comb \rfile[29][3]~feeder (
// Equation(s):
// \rfile[29][3]~feeder_combout  = \wdat_WB[3]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_3),
	.cin(gnd),
	.combout(\rfile[29][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[29][3]~feeder .lut_mask = 16'hFF00;
defparam \rfile[29][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N25
dffeas \rfile[29][3] (
	.clk(!CLK),
	.d(\rfile[29][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[29][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[29][3] .is_wysiwyg = "true";
defparam \rfile[29][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N1
dffeas \rfile[25][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][3] .is_wysiwyg = "true";
defparam \rfile[25][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N2
cycloneive_lcell_comb \rfile[17][3]~feeder (
// Equation(s):
// \rfile[17][3]~feeder_combout  = \wdat_WB[3]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[17][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[17][3]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[17][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y28_N3
dffeas \rfile[17][3] (
	.clk(!CLK),
	.d(\rfile[17][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][3] .is_wysiwyg = "true";
defparam \rfile[17][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N0
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[25][3]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[17][3]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[25][3]~q ),
	.datad(\rfile[17][3]~q ),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hB9A8;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N4
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (instruction_D[23] & ((\Mux28~0_combout  & ((\rfile[29][3]~q ))) # (!\Mux28~0_combout  & (\rfile[21][3]~q )))) # (!instruction_D[23] & (((\Mux28~0_combout ))))

	.dataa(\rfile[21][3]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[29][3]~q ),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hF388;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y36_N17
dffeas \rfile[30][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][3] .is_wysiwyg = "true";
defparam \rfile[30][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y36_N27
dffeas \rfile[22][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][3] .is_wysiwyg = "true";
defparam \rfile[22][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N20
cycloneive_lcell_comb \rfile[18][3]~feeder (
// Equation(s):
// \rfile[18][3]~feeder_combout  = \wdat_WB[3]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[18][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[18][3]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[18][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N21
dffeas \rfile[18][3] (
	.clk(!CLK),
	.d(\rfile[18][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][3] .is_wysiwyg = "true";
defparam \rfile[18][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N26
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[22][3]~q )) # (!instruction_D[23] & ((\rfile[18][3]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[22][3]~q ),
	.datad(\rfile[18][3]~q ),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hD9C8;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y36_N7
dffeas \rfile[26][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][3] .is_wysiwyg = "true";
defparam \rfile[26][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N30
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (instruction_D[24] & ((\Mux28~2_combout  & (\rfile[30][3]~q )) # (!\Mux28~2_combout  & ((\rfile[26][3]~q ))))) # (!instruction_D[24] & (((\Mux28~2_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[30][3]~q ),
	.datac(\Mux28~2_combout ),
	.datad(\rfile[26][3]~q ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hDAD0;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y32_N31
dffeas \rfile[16][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][3] .is_wysiwyg = "true";
defparam \rfile[16][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N16
cycloneive_lcell_comb \rfile[20][3]~feeder (
// Equation(s):
// \rfile[20][3]~feeder_combout  = \wdat_WB[3]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[20][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[20][3]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[20][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N17
dffeas \rfile[20][3] (
	.clk(!CLK),
	.d(\rfile[20][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][3] .is_wysiwyg = "true";
defparam \rfile[20][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N30
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[20][3]~q ))) # (!instruction_D[23] & (\rfile[16][3]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[16][3]~q ),
	.datad(\rfile[20][3]~q ),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hDC98;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y32_N29
dffeas \rfile[24][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][3] .is_wysiwyg = "true";
defparam \rfile[24][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N10
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (instruction_D[24] & ((\Mux28~4_combout  & (\rfile[28][3]~q )) # (!\Mux28~4_combout  & ((\rfile[24][3]~q ))))) # (!instruction_D[24] & (((\Mux28~4_combout ))))

	.dataa(\rfile[28][3]~q ),
	.datab(instruction_D_24),
	.datac(\Mux28~4_combout ),
	.datad(\rfile[24][3]~q ),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hBCB0;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N16
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// \Mux28~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux28~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & ((\Mux28~5_combout ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux28~3_combout ),
	.datad(\Mux28~5_combout ),
	.cin(gnd),
	.combout(\Mux28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'hB9A8;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N13
dffeas \rfile[14][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[14][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[14][3] .is_wysiwyg = "true";
defparam \rfile[14][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N5
dffeas \rfile[12][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][3] .is_wysiwyg = "true";
defparam \rfile[12][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N27
dffeas \rfile[13][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[13][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[13][3] .is_wysiwyg = "true";
defparam \rfile[13][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N4
cycloneive_lcell_comb \Mux28~17 (
// Equation(s):
// \Mux28~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][3]~q ))) # (!instruction_D[21] & (\rfile[12][3]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][3]~q ),
	.datad(\rfile[13][3]~q ),
	.cin(gnd),
	.combout(\Mux28~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~17 .lut_mask = 16'hDC98;
defparam \Mux28~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N14
cycloneive_lcell_comb \rfile[15][3]~feeder (
// Equation(s):
// \rfile[15][3]~feeder_combout  = \wdat_WB[3]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_3),
	.cin(gnd),
	.combout(\rfile[15][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[15][3]~feeder .lut_mask = 16'hFF00;
defparam \rfile[15][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N15
dffeas \rfile[15][3] (
	.clk(!CLK),
	.d(\rfile[15][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[15][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[15][3] .is_wysiwyg = "true";
defparam \rfile[15][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N24
cycloneive_lcell_comb \Mux28~18 (
// Equation(s):
// \Mux28~18_combout  = (\Mux28~17_combout  & (((\rfile[15][3]~q ) # (!instruction_D[22])))) # (!\Mux28~17_combout  & (\rfile[14][3]~q  & (instruction_D[22])))

	.dataa(\rfile[14][3]~q ),
	.datab(\Mux28~17_combout ),
	.datac(instruction_D_22),
	.datad(\rfile[15][3]~q ),
	.cin(gnd),
	.combout(\Mux28~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~18 .lut_mask = 16'hEC2C;
defparam \Mux28~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N7
dffeas \rfile[7][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][3] .is_wysiwyg = "true";
defparam \rfile[7][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N3
dffeas \rfile[4][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][3] .is_wysiwyg = "true";
defparam \rfile[4][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y28_N9
dffeas \rfile[5][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][3] .is_wysiwyg = "true";
defparam \rfile[5][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N2
cycloneive_lcell_comb \Mux28~10 (
// Equation(s):
// \Mux28~10_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[5][3]~q ))) # (!instruction_D[21] & (\rfile[4][3]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[4][3]~q ),
	.datad(\rfile[5][3]~q ),
	.cin(gnd),
	.combout(\Mux28~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~10 .lut_mask = 16'hDC98;
defparam \Mux28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N13
dffeas \rfile[6][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][3] .is_wysiwyg = "true";
defparam \rfile[6][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N12
cycloneive_lcell_comb \Mux28~11 (
// Equation(s):
// \Mux28~11_combout  = (\Mux28~10_combout  & ((\rfile[7][3]~q ) # ((!instruction_D[22])))) # (!\Mux28~10_combout  & (((\rfile[6][3]~q  & instruction_D[22]))))

	.dataa(\rfile[7][3]~q ),
	.datab(\Mux28~10_combout ),
	.datac(\rfile[6][3]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux28~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~11 .lut_mask = 16'hB8CC;
defparam \Mux28~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N1
dffeas \rfile[3][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[3][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[3][3] .is_wysiwyg = "true";
defparam \rfile[3][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N6
cycloneive_lcell_comb \rfile[1][3]~feeder (
// Equation(s):
// \rfile[1][3]~feeder_combout  = \wdat_WB[3]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_3),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[1][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[1][3]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[1][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N7
dffeas \rfile[1][3] (
	.clk(!CLK),
	.d(\rfile[1][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][3] .is_wysiwyg = "true";
defparam \rfile[1][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N0
cycloneive_lcell_comb \Mux28~14 (
// Equation(s):
// \Mux28~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][3]~q )) # (!instruction_D[22] & ((\rfile[1][3]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[3][3]~q ),
	.datad(\rfile[1][3]~q ),
	.cin(gnd),
	.combout(\Mux28~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~14 .lut_mask = 16'hC480;
defparam \Mux28~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N5
dffeas \rfile[2][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][3] .is_wysiwyg = "true";
defparam \rfile[2][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N4
cycloneive_lcell_comb \Mux28~15 (
// Equation(s):
// \Mux28~15_combout  = (\Mux28~14_combout ) # ((instruction_D[22] & (\rfile[2][3]~q  & !instruction_D[21])))

	.dataa(instruction_D_22),
	.datab(\Mux28~14_combout ),
	.datac(\rfile[2][3]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux28~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~15 .lut_mask = 16'hCCEC;
defparam \Mux28~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N25
dffeas \rfile[11][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][3] .is_wysiwyg = "true";
defparam \rfile[11][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N22
cycloneive_lcell_comb \rfile[9][3]~feeder (
// Equation(s):
// \rfile[9][3]~feeder_combout  = \wdat_WB[3]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_3),
	.cin(gnd),
	.combout(\rfile[9][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[9][3]~feeder .lut_mask = 16'hFF00;
defparam \rfile[9][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N23
dffeas \rfile[9][3] (
	.clk(!CLK),
	.d(\rfile[9][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[9][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[9][3] .is_wysiwyg = "true";
defparam \rfile[9][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N21
dffeas \rfile[10][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][3] .is_wysiwyg = "true";
defparam \rfile[10][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N20
cycloneive_lcell_comb \Mux28~12 (
// Equation(s):
// \Mux28~12_combout  = (instruction_D[21] & (((instruction_D[22])))) # (!instruction_D[21] & ((instruction_D[22] & ((\rfile[10][3]~q ))) # (!instruction_D[22] & (\rfile[8][3]~q ))))

	.dataa(\rfile[8][3]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[10][3]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux28~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~12 .lut_mask = 16'hFC22;
defparam \Mux28~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N2
cycloneive_lcell_comb \Mux28~13 (
// Equation(s):
// \Mux28~13_combout  = (instruction_D[21] & ((\Mux28~12_combout  & (\rfile[11][3]~q )) # (!\Mux28~12_combout  & ((\rfile[9][3]~q ))))) # (!instruction_D[21] & (((\Mux28~12_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[11][3]~q ),
	.datac(\rfile[9][3]~q ),
	.datad(\Mux28~12_combout ),
	.cin(gnd),
	.combout(\Mux28~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~13 .lut_mask = 16'hDDA0;
defparam \Mux28~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N18
cycloneive_lcell_comb \Mux28~16 (
// Equation(s):
// \Mux28~16_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\Mux28~13_combout )))) # (!instruction_D[24] & (!instruction_D[23] & (\Mux28~15_combout )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux28~15_combout ),
	.datad(\Mux28~13_combout ),
	.cin(gnd),
	.combout(\Mux28~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~16 .lut_mask = 16'hBA98;
defparam \Mux28~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N20
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[25][2]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[17][2]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[25][2]~q ),
	.datad(\rfile[17][2]~q ),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hB9A8;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N6
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (\Mux61~0_combout  & (((\rfile[29][2]~q ) # (!instruction_D[18])))) # (!\Mux61~0_combout  & (\rfile[21][2]~q  & ((instruction_D[18]))))

	.dataa(\rfile[21][2]~q ),
	.datab(\rfile[29][2]~q ),
	.datac(\Mux61~0_combout ),
	.datad(instruction_D_18),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hCAF0;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N12
cycloneive_lcell_comb \Mux61~7 (
// Equation(s):
// \Mux61~7_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[27][2]~q )))) # (!instruction_D[19] & (!instruction_D[18] & ((\rfile[19][2]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[27][2]~q ),
	.datad(\rfile[19][2]~q ),
	.cin(gnd),
	.combout(\Mux61~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~7 .lut_mask = 16'hB9A8;
defparam \Mux61~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N18
cycloneive_lcell_comb \Mux61~8 (
// Equation(s):
// \Mux61~8_combout  = (instruction_D[18] & ((\Mux61~7_combout  & (\rfile[31][2]~q )) # (!\Mux61~7_combout  & ((\rfile[23][2]~q ))))) # (!instruction_D[18] & (((\Mux61~7_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[31][2]~q ),
	.datac(\rfile[23][2]~q ),
	.datad(\Mux61~7_combout ),
	.cin(gnd),
	.combout(\Mux61~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~8 .lut_mask = 16'hDDA0;
defparam \Mux61~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N8
cycloneive_lcell_comb \Mux61~4 (
// Equation(s):
// \Mux61~4_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[20][2]~q )) # (!instruction_D[18] & ((\rfile[16][2]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[20][2]~q ),
	.datad(\rfile[16][2]~q ),
	.cin(gnd),
	.combout(\Mux61~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~4 .lut_mask = 16'hD9C8;
defparam \Mux61~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y32_N22
cycloneive_lcell_comb \rfile[28][2]~feeder (
// Equation(s):
// \rfile[28][2]~feeder_combout  = \wdat_WB[2]~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_2),
	.cin(gnd),
	.combout(\rfile[28][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][2]~feeder .lut_mask = 16'hFF00;
defparam \rfile[28][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X77_Y32_N23
dffeas \rfile[28][2] (
	.clk(!CLK),
	.d(\rfile[28][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][2] .is_wysiwyg = "true";
defparam \rfile[28][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N14
cycloneive_lcell_comb \Mux61~5 (
// Equation(s):
// \Mux61~5_combout  = (instruction_D[19] & ((\Mux61~4_combout  & ((\rfile[28][2]~q ))) # (!\Mux61~4_combout  & (\rfile[24][2]~q )))) # (!instruction_D[19] & (((\Mux61~4_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[24][2]~q ),
	.datac(\Mux61~4_combout ),
	.datad(\rfile[28][2]~q ),
	.cin(gnd),
	.combout(\Mux61~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~5 .lut_mask = 16'hF858;
defparam \Mux61~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y36_N22
cycloneive_lcell_comb \Mux61~2 (
// Equation(s):
// \Mux61~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[22][2]~q ))) # (!instruction_D[18] & (\rfile[18][2]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][2]~q ),
	.datad(\rfile[22][2]~q ),
	.cin(gnd),
	.combout(\Mux61~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~2 .lut_mask = 16'hDC98;
defparam \Mux61~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N24
cycloneive_lcell_comb \Mux61~3 (
// Equation(s):
// \Mux61~3_combout  = (instruction_D[19] & ((\Mux61~2_combout  & ((\rfile[30][2]~q ))) # (!\Mux61~2_combout  & (\rfile[26][2]~q )))) # (!instruction_D[19] & (((\Mux61~2_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[26][2]~q ),
	.datac(\rfile[30][2]~q ),
	.datad(\Mux61~2_combout ),
	.cin(gnd),
	.combout(\Mux61~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~3 .lut_mask = 16'hF588;
defparam \Mux61~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N20
cycloneive_lcell_comb \Mux61~6 (
// Equation(s):
// \Mux61~6_combout  = (instruction_D[17] & ((instruction_D[16]) # ((\Mux61~3_combout )))) # (!instruction_D[17] & (!instruction_D[16] & (\Mux61~5_combout )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\Mux61~5_combout ),
	.datad(\Mux61~3_combout ),
	.cin(gnd),
	.combout(\Mux61~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~6 .lut_mask = 16'hBA98;
defparam \Mux61~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N0
cycloneive_lcell_comb \Mux61~12 (
// Equation(s):
// \Mux61~12_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][2]~q ))) # (!instruction_D[17] & (\rfile[8][2]~q ))))

	.dataa(\rfile[8][2]~q ),
	.datab(instruction_D_16),
	.datac(instruction_D_17),
	.datad(\rfile[10][2]~q ),
	.cin(gnd),
	.combout(\Mux61~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~12 .lut_mask = 16'hF2C2;
defparam \Mux61~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N14
cycloneive_lcell_comb \Mux61~13 (
// Equation(s):
// \Mux61~13_combout  = (instruction_D[16] & ((\Mux61~12_combout  & (\rfile[11][2]~q )) # (!\Mux61~12_combout  & ((\rfile[9][2]~q ))))) # (!instruction_D[16] & (((\Mux61~12_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][2]~q ),
	.datac(\rfile[9][2]~q ),
	.datad(\Mux61~12_combout ),
	.cin(gnd),
	.combout(\Mux61~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~13 .lut_mask = 16'hDDA0;
defparam \Mux61~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N14
cycloneive_lcell_comb \Mux61~14 (
// Equation(s):
// \Mux61~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][2]~q ))) # (!instruction_D[17] & (\rfile[1][2]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[1][2]~q ),
	.datad(\rfile[3][2]~q ),
	.cin(gnd),
	.combout(\Mux61~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~14 .lut_mask = 16'hC840;
defparam \Mux61~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N28
cycloneive_lcell_comb \Mux61~15 (
// Equation(s):
// \Mux61~15_combout  = (\Mux61~14_combout ) # ((instruction_D[17] & (!instruction_D[16] & \rfile[2][2]~q )))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[2][2]~q ),
	.datad(\Mux61~14_combout ),
	.cin(gnd),
	.combout(\Mux61~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~15 .lut_mask = 16'hFF20;
defparam \Mux61~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N26
cycloneive_lcell_comb \Mux61~16 (
// Equation(s):
// \Mux61~16_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\Mux61~13_combout )))) # (!instruction_D[19] & (!instruction_D[18] & ((\Mux61~15_combout ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\Mux61~13_combout ),
	.datad(\Mux61~15_combout ),
	.cin(gnd),
	.combout(\Mux61~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~16 .lut_mask = 16'hB9A8;
defparam \Mux61~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N10
cycloneive_lcell_comb \Mux61~10 (
// Equation(s):
// \Mux61~10_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][2]~q ))) # (!instruction_D[16] & (\rfile[4][2]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][2]~q ),
	.datad(\rfile[5][2]~q ),
	.cin(gnd),
	.combout(\Mux61~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~10 .lut_mask = 16'hDC98;
defparam \Mux61~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N16
cycloneive_lcell_comb \Mux61~11 (
// Equation(s):
// \Mux61~11_combout  = (instruction_D[17] & ((\Mux61~10_combout  & (\rfile[7][2]~q )) # (!\Mux61~10_combout  & ((\rfile[6][2]~q ))))) # (!instruction_D[17] & (((\Mux61~10_combout ))))

	.dataa(\rfile[7][2]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[6][2]~q ),
	.datad(\Mux61~10_combout ),
	.cin(gnd),
	.combout(\Mux61~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~11 .lut_mask = 16'hBBC0;
defparam \Mux61~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N10
cycloneive_lcell_comb \Mux61~17 (
// Equation(s):
// \Mux61~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][2]~q )))) # (!instruction_D[16] & (!instruction_D[17] & ((\rfile[12][2]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[13][2]~q ),
	.datad(\rfile[12][2]~q ),
	.cin(gnd),
	.combout(\Mux61~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~17 .lut_mask = 16'hB9A8;
defparam \Mux61~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N0
cycloneive_lcell_comb \Mux61~18 (
// Equation(s):
// \Mux61~18_combout  = (instruction_D[17] & ((\Mux61~17_combout  & (\rfile[15][2]~q )) # (!\Mux61~17_combout  & ((\rfile[14][2]~q ))))) # (!instruction_D[17] & (((\Mux61~17_combout ))))

	.dataa(\rfile[15][2]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[14][2]~q ),
	.datad(\Mux61~17_combout ),
	.cin(gnd),
	.combout(\Mux61~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~18 .lut_mask = 16'hBBC0;
defparam \Mux61~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N6
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[25][8]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[17][8]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[17][8]~q ),
	.datad(\rfile[25][8]~q ),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hBA98;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N26
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (\Mux23~0_combout  & (((\rfile[29][8]~q )) # (!instruction_D[23]))) # (!\Mux23~0_combout  & (instruction_D[23] & ((\rfile[21][8]~q ))))

	.dataa(\Mux23~0_combout ),
	.datab(instruction_D_23),
	.datac(\rfile[29][8]~q ),
	.datad(\rfile[21][8]~q ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hE6A2;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N18
cycloneive_lcell_comb \Mux23~7 (
// Equation(s):
// \Mux23~7_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[27][8]~q )) # (!instruction_D[24] & ((\rfile[19][8]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[27][8]~q ),
	.datad(\rfile[19][8]~q ),
	.cin(gnd),
	.combout(\Mux23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~7 .lut_mask = 16'hD9C8;
defparam \Mux23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N22
cycloneive_lcell_comb \Mux23~8 (
// Equation(s):
// \Mux23~8_combout  = (instruction_D[23] & ((\Mux23~7_combout  & ((\rfile[31][8]~q ))) # (!\Mux23~7_combout  & (\rfile[23][8]~q )))) # (!instruction_D[23] & (((\Mux23~7_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[23][8]~q ),
	.datac(\rfile[31][8]~q ),
	.datad(\Mux23~7_combout ),
	.cin(gnd),
	.combout(\Mux23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~8 .lut_mask = 16'hF588;
defparam \Mux23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y35_N23
dffeas \rfile[30][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][8] .is_wysiwyg = "true";
defparam \rfile[30][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N18
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[22][8]~q )) # (!instruction_D[23] & ((\rfile[18][8]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[22][8]~q ),
	.datad(\rfile[18][8]~q ),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'hD9C8;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N22
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (instruction_D[24] & ((\Mux23~2_combout  & ((\rfile[30][8]~q ))) # (!\Mux23~2_combout  & (\rfile[26][8]~q )))) # (!instruction_D[24] & (((\Mux23~2_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[26][8]~q ),
	.datac(\rfile[30][8]~q ),
	.datad(\Mux23~2_combout ),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'hF588;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y30_N30
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[20][8]~q )))) # (!instruction_D[23] & (!instruction_D[24] & (\rfile[16][8]~q )))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[16][8]~q ),
	.datad(\rfile[20][8]~q ),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hBA98;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N2
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// \Mux23~5_combout  = (instruction_D[24] & ((\Mux23~4_combout  & (\rfile[28][8]~q )) # (!\Mux23~4_combout  & ((\rfile[24][8]~q ))))) # (!instruction_D[24] & (((\Mux23~4_combout ))))

	.dataa(\rfile[28][8]~q ),
	.datab(\rfile[24][8]~q ),
	.datac(instruction_D_24),
	.datad(\Mux23~4_combout ),
	.cin(gnd),
	.combout(\Mux23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hAFC0;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N28
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (instruction_D[21] & (((instruction_D[22])))) # (!instruction_D[21] & ((instruction_D[22] & (\Mux23~3_combout )) # (!instruction_D[22] & ((\Mux23~5_combout )))))

	.dataa(instruction_D_21),
	.datab(\Mux23~3_combout ),
	.datac(instruction_D_22),
	.datad(\Mux23~5_combout ),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hE5E0;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N4
cycloneive_lcell_comb \Mux23~10 (
// Equation(s):
// \Mux23~10_combout  = (instruction_D[21] & (((\rfile[5][8]~q ) # (instruction_D[22])))) # (!instruction_D[21] & (\rfile[4][8]~q  & ((!instruction_D[22]))))

	.dataa(\rfile[4][8]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[5][8]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux23~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~10 .lut_mask = 16'hCCE2;
defparam \Mux23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N8
cycloneive_lcell_comb \Mux23~11 (
// Equation(s):
// \Mux23~11_combout  = (instruction_D[22] & ((\Mux23~10_combout  & ((\rfile[7][8]~q ))) # (!\Mux23~10_combout  & (\rfile[6][8]~q )))) # (!instruction_D[22] & (((\Mux23~10_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[6][8]~q ),
	.datac(\Mux23~10_combout ),
	.datad(\rfile[7][8]~q ),
	.cin(gnd),
	.combout(\Mux23~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~11 .lut_mask = 16'hF858;
defparam \Mux23~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N8
cycloneive_lcell_comb \Mux23~12 (
// Equation(s):
// \Mux23~12_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][8]~q )))) # (!instruction_D[22] & (!instruction_D[21] & ((\rfile[8][8]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[10][8]~q ),
	.datad(\rfile[8][8]~q ),
	.cin(gnd),
	.combout(\Mux23~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~12 .lut_mask = 16'hB9A8;
defparam \Mux23~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N28
cycloneive_lcell_comb \Mux23~13 (
// Equation(s):
// \Mux23~13_combout  = (instruction_D[21] & ((\Mux23~12_combout  & ((\rfile[11][8]~q ))) # (!\Mux23~12_combout  & (\rfile[9][8]~q )))) # (!instruction_D[21] & (((\Mux23~12_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[9][8]~q ),
	.datac(\rfile[11][8]~q ),
	.datad(\Mux23~12_combout ),
	.cin(gnd),
	.combout(\Mux23~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~13 .lut_mask = 16'hF588;
defparam \Mux23~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N10
cycloneive_lcell_comb \Mux23~14 (
// Equation(s):
// \Mux23~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][8]~q ))) # (!instruction_D[22] & (\rfile[1][8]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][8]~q ),
	.datad(\rfile[3][8]~q ),
	.cin(gnd),
	.combout(\Mux23~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~14 .lut_mask = 16'hC840;
defparam \Mux23~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N20
cycloneive_lcell_comb \Mux23~15 (
// Equation(s):
// \Mux23~15_combout  = (\Mux23~14_combout ) # ((instruction_D[22] & (\rfile[2][8]~q  & !instruction_D[21])))

	.dataa(instruction_D_22),
	.datab(\rfile[2][8]~q ),
	.datac(\Mux23~14_combout ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux23~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~15 .lut_mask = 16'hF0F8;
defparam \Mux23~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N30
cycloneive_lcell_comb \Mux23~16 (
// Equation(s):
// \Mux23~16_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\Mux23~13_combout )))) # (!instruction_D[24] & (!instruction_D[23] & ((\Mux23~15_combout ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux23~13_combout ),
	.datad(\Mux23~15_combout ),
	.cin(gnd),
	.combout(\Mux23~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~16 .lut_mask = 16'hB9A8;
defparam \Mux23~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N26
cycloneive_lcell_comb \Mux23~17 (
// Equation(s):
// \Mux23~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][8]~q )) # (!instruction_D[21] & ((\rfile[12][8]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[13][8]~q ),
	.datad(\rfile[12][8]~q ),
	.cin(gnd),
	.combout(\Mux23~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~17 .lut_mask = 16'hD9C8;
defparam \Mux23~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N16
cycloneive_lcell_comb \Mux23~18 (
// Equation(s):
// \Mux23~18_combout  = (instruction_D[22] & ((\Mux23~17_combout  & ((\rfile[15][8]~q ))) # (!\Mux23~17_combout  & (\rfile[14][8]~q )))) # (!instruction_D[22] & (((\Mux23~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[14][8]~q ),
	.datac(\Mux23~17_combout ),
	.datad(\rfile[15][8]~q ),
	.cin(gnd),
	.combout(\Mux23~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~18 .lut_mask = 16'hF858;
defparam \Mux23~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N8
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (instruction_D[23] & (((\rfile[21][7]~q ) # (instruction_D[24])))) # (!instruction_D[23] & (\rfile[17][7]~q  & ((!instruction_D[24]))))

	.dataa(\rfile[17][7]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[21][7]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hCCE2;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N16
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (instruction_D[24] & ((\Mux24~0_combout  & (\rfile[29][7]~q )) # (!\Mux24~0_combout  & ((\rfile[25][7]~q ))))) # (!instruction_D[24] & (((\Mux24~0_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[29][7]~q ),
	.datac(\rfile[25][7]~q ),
	.datad(\Mux24~0_combout ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hDDA0;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N16
cycloneive_lcell_comb \Mux24~7 (
// Equation(s):
// \Mux24~7_combout  = (instruction_D[24] & (((instruction_D[23])))) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[23][7]~q ))) # (!instruction_D[23] & (\rfile[19][7]~q ))))

	.dataa(instruction_D_24),
	.datab(\rfile[19][7]~q ),
	.datac(\rfile[23][7]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~7 .lut_mask = 16'hFA44;
defparam \Mux24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N24
cycloneive_lcell_comb \Mux24~8 (
// Equation(s):
// \Mux24~8_combout  = (instruction_D[24] & ((\Mux24~7_combout  & ((\rfile[31][7]~q ))) # (!\Mux24~7_combout  & (\rfile[27][7]~q )))) # (!instruction_D[24] & (((\Mux24~7_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[27][7]~q ),
	.datac(\rfile[31][7]~q ),
	.datad(\Mux24~7_combout ),
	.cin(gnd),
	.combout(\Mux24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~8 .lut_mask = 16'hF588;
defparam \Mux24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N28
cycloneive_lcell_comb \Mux24~2 (
// Equation(s):
// \Mux24~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][7]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[18][7]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[26][7]~q ),
	.datad(\rfile[18][7]~q ),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~2 .lut_mask = 16'hB9A8;
defparam \Mux24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N20
cycloneive_lcell_comb \Mux24~3 (
// Equation(s):
// \Mux24~3_combout  = (instruction_D[23] & ((\Mux24~2_combout  & (\rfile[30][7]~q )) # (!\Mux24~2_combout  & ((\rfile[22][7]~q ))))) # (!instruction_D[23] & (((\Mux24~2_combout ))))

	.dataa(\rfile[30][7]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[22][7]~q ),
	.datad(\Mux24~2_combout ),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~3 .lut_mask = 16'hBBC0;
defparam \Mux24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N20
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (\Mux24~4_combout  & (((\rfile[28][7]~q )) # (!instruction_D[23]))) # (!\Mux24~4_combout  & (instruction_D[23] & ((\rfile[20][7]~q ))))

	.dataa(\Mux24~4_combout ),
	.datab(instruction_D_23),
	.datac(\rfile[28][7]~q ),
	.datad(\rfile[20][7]~q ),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hE6A2;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N6
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// \Mux24~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\Mux24~3_combout )) # (!instruction_D[22] & ((\Mux24~5_combout )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux24~3_combout ),
	.datad(\Mux24~5_combout ),
	.cin(gnd),
	.combout(\Mux24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'hD9C8;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N27
dffeas \rfile[12][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][7] .is_wysiwyg = "true";
defparam \rfile[12][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N26
cycloneive_lcell_comb \Mux24~17 (
// Equation(s):
// \Mux24~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][7]~q ))) # (!instruction_D[21] & (\rfile[12][7]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][7]~q ),
	.datad(\rfile[13][7]~q ),
	.cin(gnd),
	.combout(\Mux24~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~17 .lut_mask = 16'hDC98;
defparam \Mux24~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N4
cycloneive_lcell_comb \Mux24~18 (
// Equation(s):
// \Mux24~18_combout  = (instruction_D[22] & ((\Mux24~17_combout  & (\rfile[15][7]~q )) # (!\Mux24~17_combout  & ((\rfile[14][7]~q ))))) # (!instruction_D[22] & (((\Mux24~17_combout ))))

	.dataa(\rfile[15][7]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[14][7]~q ),
	.datad(\Mux24~17_combout ),
	.cin(gnd),
	.combout(\Mux24~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~18 .lut_mask = 16'hBBC0;
defparam \Mux24~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N18
cycloneive_lcell_comb \Mux24~10 (
// Equation(s):
// \Mux24~10_combout  = (instruction_D[22] & ((\rfile[10][7]~q ) # ((instruction_D[21])))) # (!instruction_D[22] & (((\rfile[8][7]~q  & !instruction_D[21]))))

	.dataa(instruction_D_22),
	.datab(\rfile[10][7]~q ),
	.datac(\rfile[8][7]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~10 .lut_mask = 16'hAAD8;
defparam \Mux24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N8
cycloneive_lcell_comb \Mux24~11 (
// Equation(s):
// \Mux24~11_combout  = (instruction_D[21] & ((\Mux24~10_combout  & ((\rfile[11][7]~q ))) # (!\Mux24~10_combout  & (\rfile[9][7]~q )))) # (!instruction_D[21] & (((\Mux24~10_combout ))))

	.dataa(\rfile[9][7]~q ),
	.datab(\rfile[11][7]~q ),
	.datac(instruction_D_21),
	.datad(\Mux24~10_combout ),
	.cin(gnd),
	.combout(\Mux24~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~11 .lut_mask = 16'hCFA0;
defparam \Mux24~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N6
cycloneive_lcell_comb \Mux24~14 (
// Equation(s):
// \Mux24~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][7]~q ))) # (!instruction_D[22] & (\rfile[1][7]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][7]~q ),
	.datad(\rfile[3][7]~q ),
	.cin(gnd),
	.combout(\Mux24~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~14 .lut_mask = 16'hC840;
defparam \Mux24~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N2
cycloneive_lcell_comb \rfile[2][7]~feeder (
// Equation(s):
// \rfile[2][7]~feeder_combout  = \wdat_WB[7]~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_7),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[2][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[2][7]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[2][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N3
dffeas \rfile[2][7] (
	.clk(!CLK),
	.d(\rfile[2][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[2][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[2][7] .is_wysiwyg = "true";
defparam \rfile[2][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N22
cycloneive_lcell_comb \Mux24~15 (
// Equation(s):
// \Mux24~15_combout  = (\Mux24~14_combout ) # ((instruction_D[22] & (\rfile[2][7]~q  & !instruction_D[21])))

	.dataa(instruction_D_22),
	.datab(\Mux24~14_combout ),
	.datac(\rfile[2][7]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux24~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~15 .lut_mask = 16'hCCEC;
defparam \Mux24~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N20
cycloneive_lcell_comb \Mux24~12 (
// Equation(s):
// \Mux24~12_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[5][7]~q ))) # (!instruction_D[21] & (\rfile[4][7]~q ))))

	.dataa(instruction_D_22),
	.datab(\rfile[4][7]~q ),
	.datac(\rfile[5][7]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux24~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~12 .lut_mask = 16'hFA44;
defparam \Mux24~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N16
cycloneive_lcell_comb \Mux24~13 (
// Equation(s):
// \Mux24~13_combout  = (instruction_D[22] & ((\Mux24~12_combout  & ((\rfile[7][7]~q ))) # (!\Mux24~12_combout  & (\rfile[6][7]~q )))) # (!instruction_D[22] & (((\Mux24~12_combout ))))

	.dataa(\rfile[6][7]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[7][7]~q ),
	.datad(\Mux24~12_combout ),
	.cin(gnd),
	.combout(\Mux24~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~13 .lut_mask = 16'hF388;
defparam \Mux24~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N10
cycloneive_lcell_comb \Mux24~16 (
// Equation(s):
// \Mux24~16_combout  = (instruction_D[23] & (((instruction_D[24]) # (\Mux24~13_combout )))) # (!instruction_D[23] & (\Mux24~15_combout  & (!instruction_D[24])))

	.dataa(instruction_D_23),
	.datab(\Mux24~15_combout ),
	.datac(instruction_D_24),
	.datad(\Mux24~13_combout ),
	.cin(gnd),
	.combout(\Mux24~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~16 .lut_mask = 16'hAEA4;
defparam \Mux24~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N4
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (instruction_D[23] & (((instruction_D[24])))) # (!instruction_D[23] & ((instruction_D[24] & ((\rfile[25][6]~q ))) # (!instruction_D[24] & (\rfile[17][6]~q ))))

	.dataa(\rfile[17][6]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[25][6]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hFC22;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N4
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\Mux25~0_combout  & ((\rfile[29][6]~q ) # ((!instruction_D[23])))) # (!\Mux25~0_combout  & (((\rfile[21][6]~q  & instruction_D[23]))))

	.dataa(\rfile[29][6]~q ),
	.datab(\Mux25~0_combout ),
	.datac(\rfile[21][6]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hB8CC;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N4
cycloneive_lcell_comb \Mux25~7 (
// Equation(s):
// \Mux25~7_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[27][6]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[19][6]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[19][6]~q ),
	.datad(\rfile[27][6]~q ),
	.cin(gnd),
	.combout(\Mux25~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~7 .lut_mask = 16'hBA98;
defparam \Mux25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N16
cycloneive_lcell_comb \Mux25~8 (
// Equation(s):
// \Mux25~8_combout  = (\Mux25~7_combout  & (((\rfile[31][6]~q ) # (!instruction_D[23])))) # (!\Mux25~7_combout  & (\rfile[23][6]~q  & ((instruction_D[23]))))

	.dataa(\rfile[23][6]~q ),
	.datab(\rfile[31][6]~q ),
	.datac(\Mux25~7_combout ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux25~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~8 .lut_mask = 16'hCAF0;
defparam \Mux25~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N28
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[20][6]~q ))) # (!instruction_D[23] & (\rfile[16][6]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[16][6]~q ),
	.datad(\rfile[20][6]~q ),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'hDC98;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N20
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// \Mux25~5_combout  = (instruction_D[24] & ((\Mux25~4_combout  & (\rfile[28][6]~q )) # (!\Mux25~4_combout  & ((\rfile[24][6]~q ))))) # (!instruction_D[24] & (((\Mux25~4_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[28][6]~q ),
	.datac(\rfile[24][6]~q ),
	.datad(\Mux25~4_combout ),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hDDA0;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y35_N9
dffeas \rfile[26][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][6] .is_wysiwyg = "true";
defparam \rfile[26][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N8
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (\Mux25~2_combout  & (((\rfile[30][6]~q )) # (!instruction_D[24]))) # (!\Mux25~2_combout  & (instruction_D[24] & (\rfile[26][6]~q )))

	.dataa(\Mux25~2_combout ),
	.datab(instruction_D_24),
	.datac(\rfile[26][6]~q ),
	.datad(\rfile[30][6]~q ),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'hEA62;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N24
cycloneive_lcell_comb \Mux25~6 (
// Equation(s):
// \Mux25~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & ((\Mux25~3_combout ))) # (!instruction_D[22] & (\Mux25~5_combout ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux25~5_combout ),
	.datad(\Mux25~3_combout ),
	.cin(gnd),
	.combout(\Mux25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~6 .lut_mask = 16'hDC98;
defparam \Mux25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y28_N31
dffeas \rfile[4][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][6] .is_wysiwyg = "true";
defparam \rfile[4][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N30
cycloneive_lcell_comb \Mux25~10 (
// Equation(s):
// \Mux25~10_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[5][6]~q ))) # (!instruction_D[21] & (\rfile[4][6]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[4][6]~q ),
	.datad(\rfile[5][6]~q ),
	.cin(gnd),
	.combout(\Mux25~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~10 .lut_mask = 16'hDC98;
defparam \Mux25~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N18
cycloneive_lcell_comb \Mux25~11 (
// Equation(s):
// \Mux25~11_combout  = (instruction_D[22] & ((\Mux25~10_combout  & ((\rfile[7][6]~q ))) # (!\Mux25~10_combout  & (\rfile[6][6]~q )))) # (!instruction_D[22] & (((\Mux25~10_combout ))))

	.dataa(\rfile[6][6]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[7][6]~q ),
	.datad(\Mux25~10_combout ),
	.cin(gnd),
	.combout(\Mux25~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~11 .lut_mask = 16'hF388;
defparam \Mux25~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N12
cycloneive_lcell_comb \Mux25~14 (
// Equation(s):
// \Mux25~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][6]~q ))) # (!instruction_D[22] & (\rfile[1][6]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][6]~q ),
	.datad(\rfile[3][6]~q ),
	.cin(gnd),
	.combout(\Mux25~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~14 .lut_mask = 16'hC840;
defparam \Mux25~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N26
cycloneive_lcell_comb \Mux25~15 (
// Equation(s):
// \Mux25~15_combout  = (\Mux25~14_combout ) # ((\rfile[2][6]~q  & (instruction_D[22] & !instruction_D[21])))

	.dataa(\rfile[2][6]~q ),
	.datab(instruction_D_22),
	.datac(instruction_D_21),
	.datad(\Mux25~14_combout ),
	.cin(gnd),
	.combout(\Mux25~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~15 .lut_mask = 16'hFF08;
defparam \Mux25~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N20
cycloneive_lcell_comb \rfile[11][6]~feeder (
// Equation(s):
// \rfile[11][6]~feeder_combout  = \wdat_WB[6]~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_6),
	.cin(gnd),
	.combout(\rfile[11][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[11][6]~feeder .lut_mask = 16'hFF00;
defparam \rfile[11][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y27_N21
dffeas \rfile[11][6] (
	.clk(!CLK),
	.d(\rfile[11][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][6] .is_wysiwyg = "true";
defparam \rfile[11][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N28
cycloneive_lcell_comb \Mux25~12 (
// Equation(s):
// \Mux25~12_combout  = (instruction_D[21] & (((instruction_D[22])))) # (!instruction_D[21] & ((instruction_D[22] & (\rfile[10][6]~q )) # (!instruction_D[22] & ((\rfile[8][6]~q )))))

	.dataa(\rfile[10][6]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[8][6]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux25~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~12 .lut_mask = 16'hEE30;
defparam \Mux25~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N0
cycloneive_lcell_comb \Mux25~13 (
// Equation(s):
// \Mux25~13_combout  = (instruction_D[21] & ((\Mux25~12_combout  & (\rfile[11][6]~q )) # (!\Mux25~12_combout  & ((\rfile[9][6]~q ))))) # (!instruction_D[21] & (((\Mux25~12_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[11][6]~q ),
	.datac(\Mux25~12_combout ),
	.datad(\rfile[9][6]~q ),
	.cin(gnd),
	.combout(\Mux25~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~13 .lut_mask = 16'hDAD0;
defparam \Mux25~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N4
cycloneive_lcell_comb \Mux25~16 (
// Equation(s):
// \Mux25~16_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\Mux25~13_combout ))) # (!instruction_D[24] & (\Mux25~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux25~15_combout ),
	.datad(\Mux25~13_combout ),
	.cin(gnd),
	.combout(\Mux25~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~16 .lut_mask = 16'hDC98;
defparam \Mux25~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N12
cycloneive_lcell_comb \Mux25~17 (
// Equation(s):
// \Mux25~17_combout  = (instruction_D[21] & (((\rfile[13][6]~q ) # (instruction_D[22])))) # (!instruction_D[21] & (\rfile[12][6]~q  & ((!instruction_D[22]))))

	.dataa(\rfile[12][6]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[13][6]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux25~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~17 .lut_mask = 16'hCCE2;
defparam \Mux25~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N22
cycloneive_lcell_comb \Mux25~18 (
// Equation(s):
// \Mux25~18_combout  = (instruction_D[22] & ((\Mux25~17_combout  & (\rfile[15][6]~q )) # (!\Mux25~17_combout  & ((\rfile[14][6]~q ))))) # (!instruction_D[22] & (((\Mux25~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[15][6]~q ),
	.datac(\Mux25~17_combout ),
	.datad(\rfile[14][6]~q ),
	.cin(gnd),
	.combout(\Mux25~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~18 .lut_mask = 16'hDAD0;
defparam \Mux25~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y27_N2
cycloneive_lcell_comb \Mux26~7 (
// Equation(s):
// \Mux26~7_combout  = (instruction_D[24] & (((instruction_D[23])))) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[23][5]~q ))) # (!instruction_D[23] & (\rfile[19][5]~q ))))

	.dataa(instruction_D_24),
	.datab(\rfile[19][5]~q ),
	.datac(instruction_D_23),
	.datad(\rfile[23][5]~q ),
	.cin(gnd),
	.combout(\Mux26~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~7 .lut_mask = 16'hF4A4;
defparam \Mux26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N26
cycloneive_lcell_comb \Mux26~8 (
// Equation(s):
// \Mux26~8_combout  = (instruction_D[24] & ((\Mux26~7_combout  & (\rfile[31][5]~q )) # (!\Mux26~7_combout  & ((\rfile[27][5]~q ))))) # (!instruction_D[24] & (((\Mux26~7_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[31][5]~q ),
	.datac(\rfile[27][5]~q ),
	.datad(\Mux26~7_combout ),
	.cin(gnd),
	.combout(\Mux26~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~8 .lut_mask = 16'hDDA0;
defparam \Mux26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N15
dffeas \rfile[22][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][5] .is_wysiwyg = "true";
defparam \rfile[22][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N0
cycloneive_lcell_comb \rfile[18][5]~feeder (
// Equation(s):
// \rfile[18][5]~feeder_combout  = \wdat_WB[5]~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_5),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[18][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[18][5]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[18][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N1
dffeas \rfile[18][5] (
	.clk(!CLK),
	.d(\rfile[18][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][5] .is_wysiwyg = "true";
defparam \rfile[18][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N2
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][5]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[18][5]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][5]~q ),
	.datad(\rfile[26][5]~q ),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'hBA98;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N14
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (instruction_D[23] & ((\Mux26~2_combout  & (\rfile[30][5]~q )) # (!\Mux26~2_combout  & ((\rfile[22][5]~q ))))) # (!instruction_D[23] & (((\Mux26~2_combout ))))

	.dataa(\rfile[30][5]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[22][5]~q ),
	.datad(\Mux26~2_combout ),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'hBBC0;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y32_N17
dffeas \rfile[28][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][5] .is_wysiwyg = "true";
defparam \rfile[28][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N2
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[24][5]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[16][5]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[16][5]~q ),
	.datad(\rfile[24][5]~q ),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'hBA98;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N16
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// \Mux26~5_combout  = (instruction_D[23] & ((\Mux26~4_combout  & ((\rfile[28][5]~q ))) # (!\Mux26~4_combout  & (\rfile[20][5]~q )))) # (!instruction_D[23] & (((\Mux26~4_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[20][5]~q ),
	.datac(\rfile[28][5]~q ),
	.datad(\Mux26~4_combout ),
	.cin(gnd),
	.combout(\Mux26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hF588;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N4
cycloneive_lcell_comb \Mux26~6 (
// Equation(s):
// \Mux26~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\Mux26~3_combout )) # (!instruction_D[22] & ((\Mux26~5_combout )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux26~3_combout ),
	.datad(\Mux26~5_combout ),
	.cin(gnd),
	.combout(\Mux26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~6 .lut_mask = 16'hD9C8;
defparam \Mux26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N2
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[21][5]~q )) # (!instruction_D[23] & ((\rfile[17][5]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[21][5]~q ),
	.datad(\rfile[17][5]~q ),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hD9C8;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N20
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (instruction_D[24] & ((\Mux26~0_combout  & (\rfile[29][5]~q )) # (!\Mux26~0_combout  & ((\rfile[25][5]~q ))))) # (!instruction_D[24] & (\Mux26~0_combout ))

	.dataa(instruction_D_24),
	.datab(\Mux26~0_combout ),
	.datac(\rfile[29][5]~q ),
	.datad(\rfile[25][5]~q ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hE6C4;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N18
cycloneive_lcell_comb \Mux26~12 (
// Equation(s):
// \Mux26~12_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[5][5]~q ))) # (!instruction_D[21] & (\rfile[4][5]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[4][5]~q ),
	.datad(\rfile[5][5]~q ),
	.cin(gnd),
	.combout(\Mux26~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~12 .lut_mask = 16'hDC98;
defparam \Mux26~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N4
cycloneive_lcell_comb \Mux26~13 (
// Equation(s):
// \Mux26~13_combout  = (\Mux26~12_combout  & ((\rfile[7][5]~q ) # ((!instruction_D[22])))) # (!\Mux26~12_combout  & (((\rfile[6][5]~q  & instruction_D[22]))))

	.dataa(\rfile[7][5]~q ),
	.datab(\rfile[6][5]~q ),
	.datac(\Mux26~12_combout ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux26~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~13 .lut_mask = 16'hACF0;
defparam \Mux26~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N28
cycloneive_lcell_comb \Mux26~14 (
// Equation(s):
// \Mux26~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][5]~q ))) # (!instruction_D[22] & (\rfile[1][5]~q ))))

	.dataa(\rfile[1][5]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[3][5]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux26~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~14 .lut_mask = 16'hE200;
defparam \Mux26~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N18
cycloneive_lcell_comb \Mux26~15 (
// Equation(s):
// \Mux26~15_combout  = (\Mux26~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][5]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[2][5]~q ),
	.datad(\Mux26~14_combout ),
	.cin(gnd),
	.combout(\Mux26~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~15 .lut_mask = 16'hFF20;
defparam \Mux26~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N12
cycloneive_lcell_comb \Mux26~16 (
// Equation(s):
// \Mux26~16_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\Mux26~13_combout )))) # (!instruction_D[23] & (!instruction_D[24] & ((\Mux26~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux26~13_combout ),
	.datad(\Mux26~15_combout ),
	.cin(gnd),
	.combout(\Mux26~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~16 .lut_mask = 16'hB9A8;
defparam \Mux26~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N12
cycloneive_lcell_comb \Mux26~10 (
// Equation(s):
// \Mux26~10_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][5]~q )))) # (!instruction_D[22] & (!instruction_D[21] & (\rfile[8][5]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[8][5]~q ),
	.datad(\rfile[10][5]~q ),
	.cin(gnd),
	.combout(\Mux26~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~10 .lut_mask = 16'hBA98;
defparam \Mux26~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N10
cycloneive_lcell_comb \Mux26~11 (
// Equation(s):
// \Mux26~11_combout  = (instruction_D[21] & ((\Mux26~10_combout  & ((\rfile[11][5]~q ))) # (!\Mux26~10_combout  & (\rfile[9][5]~q )))) # (!instruction_D[21] & (((\Mux26~10_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[9][5]~q ),
	.datac(\Mux26~10_combout ),
	.datad(\rfile[11][5]~q ),
	.cin(gnd),
	.combout(\Mux26~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~11 .lut_mask = 16'hF858;
defparam \Mux26~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N0
cycloneive_lcell_comb \Mux26~17 (
// Equation(s):
// \Mux26~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][5]~q ))) # (!instruction_D[21] & (\rfile[12][5]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][5]~q ),
	.datad(\rfile[13][5]~q ),
	.cin(gnd),
	.combout(\Mux26~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~17 .lut_mask = 16'hDC98;
defparam \Mux26~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N2
cycloneive_lcell_comb \Mux26~18 (
// Equation(s):
// \Mux26~18_combout  = (instruction_D[22] & ((\Mux26~17_combout  & ((\rfile[15][5]~q ))) # (!\Mux26~17_combout  & (\rfile[14][5]~q )))) # (!instruction_D[22] & (((\Mux26~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[14][5]~q ),
	.datac(\rfile[15][5]~q ),
	.datad(\Mux26~17_combout ),
	.cin(gnd),
	.combout(\Mux26~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~18 .lut_mask = 16'hF588;
defparam \Mux26~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y29_N23
dffeas \rfile[19][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][3] .is_wysiwyg = "true";
defparam \rfile[19][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N22
cycloneive_lcell_comb \Mux60~7 (
// Equation(s):
// \Mux60~7_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[23][3]~q ))) # (!instruction_D[18] & (\rfile[19][3]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[19][3]~q ),
	.datad(\rfile[23][3]~q ),
	.cin(gnd),
	.combout(\Mux60~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~7 .lut_mask = 16'hDC98;
defparam \Mux60~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N28
cycloneive_lcell_comb \Mux60~8 (
// Equation(s):
// \Mux60~8_combout  = (\Mux60~7_combout  & (((\rfile[31][3]~q )) # (!instruction_D[19]))) # (!\Mux60~7_combout  & (instruction_D[19] & (\rfile[27][3]~q )))

	.dataa(\Mux60~7_combout ),
	.datab(instruction_D_19),
	.datac(\rfile[27][3]~q ),
	.datad(\rfile[31][3]~q ),
	.cin(gnd),
	.combout(\Mux60~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~8 .lut_mask = 16'hEA62;
defparam \Mux60~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N30
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\rfile[21][3]~q )))) # (!instruction_D[18] & (!instruction_D[19] & ((\rfile[17][3]~q ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[21][3]~q ),
	.datad(\rfile[17][3]~q ),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'hB9A8;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N8
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (\Mux60~0_combout  & (((\rfile[29][3]~q ) # (!instruction_D[19])))) # (!\Mux60~0_combout  & (\rfile[25][3]~q  & (instruction_D[19])))

	.dataa(\Mux60~0_combout ),
	.datab(\rfile[25][3]~q ),
	.datac(instruction_D_19),
	.datad(\rfile[29][3]~q ),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hEA4A;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N6
cycloneive_lcell_comb \Mux60~2 (
// Equation(s):
// \Mux60~2_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[26][3]~q )) # (!instruction_D[19] & ((\rfile[18][3]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[26][3]~q ),
	.datad(\rfile[18][3]~q ),
	.cin(gnd),
	.combout(\Mux60~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~2 .lut_mask = 16'hD9C8;
defparam \Mux60~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N16
cycloneive_lcell_comb \Mux60~3 (
// Equation(s):
// \Mux60~3_combout  = (instruction_D[18] & ((\Mux60~2_combout  & ((\rfile[30][3]~q ))) # (!\Mux60~2_combout  & (\rfile[22][3]~q )))) # (!instruction_D[18] & (((\Mux60~2_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[22][3]~q ),
	.datac(\rfile[30][3]~q ),
	.datad(\Mux60~2_combout ),
	.cin(gnd),
	.combout(\Mux60~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~3 .lut_mask = 16'hF588;
defparam \Mux60~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N7
dffeas \rfile[28][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][3] .is_wysiwyg = "true";
defparam \rfile[28][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N28
cycloneive_lcell_comb \Mux60~4 (
// Equation(s):
// \Mux60~4_combout  = (instruction_D[18] & (((instruction_D[19])))) # (!instruction_D[18] & ((instruction_D[19] & ((\rfile[24][3]~q ))) # (!instruction_D[19] & (\rfile[16][3]~q ))))

	.dataa(\rfile[16][3]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[24][3]~q ),
	.datad(instruction_D_19),
	.cin(gnd),
	.combout(\Mux60~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~4 .lut_mask = 16'hFC22;
defparam \Mux60~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N6
cycloneive_lcell_comb \Mux60~5 (
// Equation(s):
// \Mux60~5_combout  = (instruction_D[18] & ((\Mux60~4_combout  & ((\rfile[28][3]~q ))) # (!\Mux60~4_combout  & (\rfile[20][3]~q )))) # (!instruction_D[18] & (((\Mux60~4_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[20][3]~q ),
	.datac(\rfile[28][3]~q ),
	.datad(\Mux60~4_combout ),
	.cin(gnd),
	.combout(\Mux60~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~5 .lut_mask = 16'hF588;
defparam \Mux60~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N6
cycloneive_lcell_comb \Mux60~6 (
// Equation(s):
// \Mux60~6_combout  = (instruction_D[17] & ((\Mux60~3_combout ) # ((instruction_D[16])))) # (!instruction_D[17] & (((!instruction_D[16] & \Mux60~5_combout ))))

	.dataa(instruction_D_17),
	.datab(\Mux60~3_combout ),
	.datac(instruction_D_16),
	.datad(\Mux60~5_combout ),
	.cin(gnd),
	.combout(\Mux60~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~6 .lut_mask = 16'hADA8;
defparam \Mux60~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N8
cycloneive_lcell_comb \Mux60~12 (
// Equation(s):
// \Mux60~12_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & (\rfile[5][3]~q )) # (!instruction_D[16] & ((\rfile[4][3]~q )))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[5][3]~q ),
	.datad(\rfile[4][3]~q ),
	.cin(gnd),
	.combout(\Mux60~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~12 .lut_mask = 16'hD9C8;
defparam \Mux60~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N6
cycloneive_lcell_comb \Mux60~13 (
// Equation(s):
// \Mux60~13_combout  = (instruction_D[17] & ((\Mux60~12_combout  & ((\rfile[7][3]~q ))) # (!\Mux60~12_combout  & (\rfile[6][3]~q )))) # (!instruction_D[17] & (((\Mux60~12_combout ))))

	.dataa(\rfile[6][3]~q ),
	.datab(instruction_D_17),
	.datac(\rfile[7][3]~q ),
	.datad(\Mux60~12_combout ),
	.cin(gnd),
	.combout(\Mux60~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~13 .lut_mask = 16'hF388;
defparam \Mux60~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N24
cycloneive_lcell_comb \Mux60~14 (
// Equation(s):
// \Mux60~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][3]~q ))) # (!instruction_D[17] & (\rfile[1][3]~q ))))

	.dataa(\rfile[1][3]~q ),
	.datab(\rfile[3][3]~q ),
	.datac(instruction_D_17),
	.datad(instruction_D_16),
	.cin(gnd),
	.combout(\Mux60~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~14 .lut_mask = 16'hCA00;
defparam \Mux60~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N0
cycloneive_lcell_comb \Mux60~15 (
// Equation(s):
// \Mux60~15_combout  = (\Mux60~14_combout ) # ((!instruction_D[16] & (\rfile[2][3]~q  & instruction_D[17])))

	.dataa(instruction_D_16),
	.datab(\rfile[2][3]~q ),
	.datac(instruction_D_17),
	.datad(\Mux60~14_combout ),
	.cin(gnd),
	.combout(\Mux60~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~15 .lut_mask = 16'hFF40;
defparam \Mux60~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N14
cycloneive_lcell_comb \Mux60~16 (
// Equation(s):
// \Mux60~16_combout  = (instruction_D[18] & ((instruction_D[19]) # ((\Mux60~13_combout )))) # (!instruction_D[18] & (!instruction_D[19] & ((\Mux60~15_combout ))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\Mux60~13_combout ),
	.datad(\Mux60~15_combout ),
	.cin(gnd),
	.combout(\Mux60~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~16 .lut_mask = 16'hB9A8;
defparam \Mux60~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N7
dffeas \rfile[8][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][3] .is_wysiwyg = "true";
defparam \rfile[8][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N6
cycloneive_lcell_comb \Mux60~10 (
// Equation(s):
// \Mux60~10_combout  = (instruction_D[16] & (((instruction_D[17])))) # (!instruction_D[16] & ((instruction_D[17] & (\rfile[10][3]~q )) # (!instruction_D[17] & ((\rfile[8][3]~q )))))

	.dataa(instruction_D_16),
	.datab(\rfile[10][3]~q ),
	.datac(\rfile[8][3]~q ),
	.datad(instruction_D_17),
	.cin(gnd),
	.combout(\Mux60~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~10 .lut_mask = 16'hEE50;
defparam \Mux60~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N0
cycloneive_lcell_comb \Mux60~11 (
// Equation(s):
// \Mux60~11_combout  = (instruction_D[16] & ((\Mux60~10_combout  & (\rfile[11][3]~q )) # (!\Mux60~10_combout  & ((\rfile[9][3]~q ))))) # (!instruction_D[16] & (((\Mux60~10_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][3]~q ),
	.datac(\Mux60~10_combout ),
	.datad(\rfile[9][3]~q ),
	.cin(gnd),
	.combout(\Mux60~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~11 .lut_mask = 16'hDAD0;
defparam \Mux60~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N26
cycloneive_lcell_comb \Mux60~17 (
// Equation(s):
// \Mux60~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][3]~q )))) # (!instruction_D[16] & (!instruction_D[17] & ((\rfile[12][3]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[13][3]~q ),
	.datad(\rfile[12][3]~q ),
	.cin(gnd),
	.combout(\Mux60~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~17 .lut_mask = 16'hB9A8;
defparam \Mux60~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N12
cycloneive_lcell_comb \Mux60~18 (
// Equation(s):
// \Mux60~18_combout  = (\Mux60~17_combout  & (((\rfile[15][3]~q )) # (!instruction_D[17]))) # (!\Mux60~17_combout  & (instruction_D[17] & (\rfile[14][3]~q )))

	.dataa(\Mux60~17_combout ),
	.datab(instruction_D_17),
	.datac(\rfile[14][3]~q ),
	.datad(\rfile[15][3]~q ),
	.cin(gnd),
	.combout(\Mux60~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~18 .lut_mask = 16'hEA62;
defparam \Mux60~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N12
cycloneive_lcell_comb \Mux15~7 (
// Equation(s):
// \Mux15~7_combout  = (instruction_D[24] & (((\rfile[27][16]~q ) # (instruction_D[23])))) # (!instruction_D[24] & (\rfile[19][16]~q  & ((!instruction_D[23]))))

	.dataa(\rfile[19][16]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[27][16]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~7 .lut_mask = 16'hCCE2;
defparam \Mux15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N6
cycloneive_lcell_comb \Mux15~8 (
// Equation(s):
// \Mux15~8_combout  = (instruction_D[23] & ((\Mux15~7_combout  & ((\rfile[31][16]~q ))) # (!\Mux15~7_combout  & (\rfile[23][16]~q )))) # (!instruction_D[23] & (((\Mux15~7_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[23][16]~q ),
	.datac(\rfile[31][16]~q ),
	.datad(\Mux15~7_combout ),
	.cin(gnd),
	.combout(\Mux15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~8 .lut_mask = 16'hF588;
defparam \Mux15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N4
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// \Mux15~4_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[20][16]~q )))) # (!instruction_D[23] & (!instruction_D[24] & ((\rfile[16][16]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[20][16]~q ),
	.datad(\rfile[16][16]~q ),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hB9A8;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N24
cycloneive_lcell_comb \Mux15~5 (
// Equation(s):
// \Mux15~5_combout  = (instruction_D[24] & ((\Mux15~4_combout  & ((\rfile[28][16]~q ))) # (!\Mux15~4_combout  & (\rfile[24][16]~q )))) # (!instruction_D[24] & (((\Mux15~4_combout ))))

	.dataa(\rfile[24][16]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[28][16]~q ),
	.datad(\Mux15~4_combout ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~5 .lut_mask = 16'hF388;
defparam \Mux15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N26
cycloneive_lcell_comb \rfile[22][16]~feeder (
// Equation(s):
// \rfile[22][16]~feeder_combout  = \wdat_WB[16]~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_16),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[22][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[22][16]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[22][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y35_N27
dffeas \rfile[22][16] (
	.clk(!CLK),
	.d(\rfile[22][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][16] .is_wysiwyg = "true";
defparam \rfile[22][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N31
dffeas \rfile[18][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][16] .is_wysiwyg = "true";
defparam \rfile[18][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N2
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[22][16]~q )) # (!instruction_D[23] & ((\rfile[18][16]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[22][16]~q ),
	.datad(\rfile[18][16]~q ),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'hD9C8;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N12
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (instruction_D[24] & ((\Mux15~2_combout  & ((\rfile[30][16]~q ))) # (!\Mux15~2_combout  & (\rfile[26][16]~q )))) # (!instruction_D[24] & (((\Mux15~2_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[26][16]~q ),
	.datac(\rfile[30][16]~q ),
	.datad(\Mux15~2_combout ),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hF588;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N14
cycloneive_lcell_comb \Mux15~6 (
// Equation(s):
// \Mux15~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & ((\Mux15~3_combout ))) # (!instruction_D[22] & (\Mux15~5_combout ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux15~5_combout ),
	.datad(\Mux15~3_combout ),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~6 .lut_mask = 16'hDC98;
defparam \Mux15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N18
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[25][16]~q )) # (!instruction_D[24] & ((\rfile[17][16]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[25][16]~q ),
	.datad(\rfile[17][16]~q ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hD9C8;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N14
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (instruction_D[23] & ((\Mux15~0_combout  & ((\rfile[29][16]~q ))) # (!\Mux15~0_combout  & (\rfile[21][16]~q )))) # (!instruction_D[23] & (((\Mux15~0_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[21][16]~q ),
	.datac(\rfile[29][16]~q ),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hF588;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y28_N27
dffeas \rfile[4][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][16] .is_wysiwyg = "true";
defparam \rfile[4][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N26
cycloneive_lcell_comb \Mux15~10 (
// Equation(s):
// \Mux15~10_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[5][16]~q ))) # (!instruction_D[21] & (\rfile[4][16]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[4][16]~q ),
	.datad(\rfile[5][16]~q ),
	.cin(gnd),
	.combout(\Mux15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~10 .lut_mask = 16'hDC98;
defparam \Mux15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N2
cycloneive_lcell_comb \Mux15~11 (
// Equation(s):
// \Mux15~11_combout  = (\Mux15~10_combout  & (((\rfile[7][16]~q ) # (!instruction_D[22])))) # (!\Mux15~10_combout  & (\rfile[6][16]~q  & ((instruction_D[22]))))

	.dataa(\rfile[6][16]~q ),
	.datab(\rfile[7][16]~q ),
	.datac(\Mux15~10_combout ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux15~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~11 .lut_mask = 16'hCAF0;
defparam \Mux15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N16
cycloneive_lcell_comb \Mux15~14 (
// Equation(s):
// \Mux15~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][16]~q ))) # (!instruction_D[22] & (\rfile[1][16]~q ))))

	.dataa(\rfile[1][16]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[3][16]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux15~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~14 .lut_mask = 16'hE200;
defparam \Mux15~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N4
cycloneive_lcell_comb \Mux15~15 (
// Equation(s):
// \Mux15~15_combout  = (\Mux15~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][16]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[2][16]~q ),
	.datad(\Mux15~14_combout ),
	.cin(gnd),
	.combout(\Mux15~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~15 .lut_mask = 16'hFF20;
defparam \Mux15~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y35_N23
dffeas \rfile[8][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][16] .is_wysiwyg = "true";
defparam \rfile[8][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N22
cycloneive_lcell_comb \Mux15~12 (
// Equation(s):
// \Mux15~12_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][16]~q )))) # (!instruction_D[22] & (!instruction_D[21] & (\rfile[8][16]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[8][16]~q ),
	.datad(\rfile[10][16]~q ),
	.cin(gnd),
	.combout(\Mux15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~12 .lut_mask = 16'hBA98;
defparam \Mux15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N2
cycloneive_lcell_comb \Mux15~13 (
// Equation(s):
// \Mux15~13_combout  = (instruction_D[21] & ((\Mux15~12_combout  & ((\rfile[11][16]~q ))) # (!\Mux15~12_combout  & (\rfile[9][16]~q )))) # (!instruction_D[21] & (((\Mux15~12_combout ))))

	.dataa(\rfile[9][16]~q ),
	.datab(\rfile[11][16]~q ),
	.datac(instruction_D_21),
	.datad(\Mux15~12_combout ),
	.cin(gnd),
	.combout(\Mux15~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~13 .lut_mask = 16'hCFA0;
defparam \Mux15~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N30
cycloneive_lcell_comb \Mux15~16 (
// Equation(s):
// \Mux15~16_combout  = (instruction_D[24] & (((instruction_D[23]) # (\Mux15~13_combout )))) # (!instruction_D[24] & (\Mux15~15_combout  & (!instruction_D[23])))

	.dataa(instruction_D_24),
	.datab(\Mux15~15_combout ),
	.datac(instruction_D_23),
	.datad(\Mux15~13_combout ),
	.cin(gnd),
	.combout(\Mux15~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~16 .lut_mask = 16'hAEA4;
defparam \Mux15~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N22
cycloneive_lcell_comb \Mux15~17 (
// Equation(s):
// \Mux15~17_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][16]~q ))) # (!instruction_D[21] & (\rfile[12][16]~q ))))

	.dataa(instruction_D_22),
	.datab(\rfile[12][16]~q ),
	.datac(instruction_D_21),
	.datad(\rfile[13][16]~q ),
	.cin(gnd),
	.combout(\Mux15~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~17 .lut_mask = 16'hF4A4;
defparam \Mux15~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N24
cycloneive_lcell_comb \Mux15~18 (
// Equation(s):
// \Mux15~18_combout  = (instruction_D[22] & ((\Mux15~17_combout  & (\rfile[15][16]~q )) # (!\Mux15~17_combout  & ((\rfile[14][16]~q ))))) # (!instruction_D[22] & (((\Mux15~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[15][16]~q ),
	.datac(\Mux15~17_combout ),
	.datad(\rfile[14][16]~q ),
	.cin(gnd),
	.combout(\Mux15~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~18 .lut_mask = 16'hDAD0;
defparam \Mux15~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N2
cycloneive_lcell_comb \Mux16~7 (
// Equation(s):
// \Mux16~7_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[23][15]~q ))) # (!instruction_D[23] & (\rfile[19][15]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[19][15]~q ),
	.datad(\rfile[23][15]~q ),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~7 .lut_mask = 16'hDC98;
defparam \Mux16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N16
cycloneive_lcell_comb \Mux16~8 (
// Equation(s):
// \Mux16~8_combout  = (instruction_D[24] & ((\Mux16~7_combout  & (\rfile[31][15]~q )) # (!\Mux16~7_combout  & ((\rfile[27][15]~q ))))) # (!instruction_D[24] & (((\Mux16~7_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[31][15]~q ),
	.datac(\rfile[27][15]~q ),
	.datad(\Mux16~7_combout ),
	.cin(gnd),
	.combout(\Mux16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~8 .lut_mask = 16'hDDA0;
defparam \Mux16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N28
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[21][15]~q )) # (!instruction_D[23] & ((\rfile[17][15]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[21][15]~q ),
	.datad(\rfile[17][15]~q ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hD9C8;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N10
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (instruction_D[24] & ((\Mux16~0_combout  & ((\rfile[29][15]~q ))) # (!\Mux16~0_combout  & (\rfile[25][15]~q )))) # (!instruction_D[24] & (((\Mux16~0_combout ))))

	.dataa(\rfile[25][15]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[29][15]~q ),
	.datad(\Mux16~0_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hF388;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N26
cycloneive_lcell_comb \rfile[28][15]~feeder (
// Equation(s):
// \rfile[28][15]~feeder_combout  = \wdat_WB[15]~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_15),
	.cin(gnd),
	.combout(\rfile[28][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][15]~feeder .lut_mask = 16'hFF00;
defparam \rfile[28][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y32_N27
dffeas \rfile[28][15] (
	.clk(!CLK),
	.d(\rfile[28][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][15] .is_wysiwyg = "true";
defparam \rfile[28][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y33_N31
dffeas \rfile[24][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][15] .is_wysiwyg = "true";
defparam \rfile[24][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N30
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[24][15]~q )) # (!instruction_D[24] & ((\rfile[16][15]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[24][15]~q ),
	.datad(\rfile[16][15]~q ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hD9C8;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N2
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// \Mux16~5_combout  = (instruction_D[23] & ((\Mux16~4_combout  & (\rfile[28][15]~q )) # (!\Mux16~4_combout  & ((\rfile[20][15]~q ))))) # (!instruction_D[23] & (((\Mux16~4_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[28][15]~q ),
	.datac(\Mux16~4_combout ),
	.datad(\rfile[20][15]~q ),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hDAD0;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N20
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[26][15]~q )) # (!instruction_D[24] & ((\rfile[18][15]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[26][15]~q ),
	.datad(\rfile[18][15]~q ),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hD9C8;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N0
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (instruction_D[23] & ((\Mux16~2_combout  & (\rfile[30][15]~q )) # (!\Mux16~2_combout  & ((\rfile[22][15]~q ))))) # (!instruction_D[23] & (((\Mux16~2_combout ))))

	.dataa(\rfile[30][15]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[22][15]~q ),
	.datad(\Mux16~2_combout ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hBBC0;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N2
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// \Mux16~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & ((\Mux16~3_combout ))) # (!instruction_D[22] & (\Mux16~5_combout ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux16~5_combout ),
	.datad(\Mux16~3_combout ),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'hDC98;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N14
cycloneive_lcell_comb \Mux16~17 (
// Equation(s):
// \Mux16~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][15]~q ))) # (!instruction_D[21] & (\rfile[12][15]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][15]~q ),
	.datad(\rfile[13][15]~q ),
	.cin(gnd),
	.combout(\Mux16~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~17 .lut_mask = 16'hDC98;
defparam \Mux16~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N2
cycloneive_lcell_comb \Mux16~18 (
// Equation(s):
// \Mux16~18_combout  = (instruction_D[22] & ((\Mux16~17_combout  & (\rfile[15][15]~q )) # (!\Mux16~17_combout  & ((\rfile[14][15]~q ))))) # (!instruction_D[22] & (((\Mux16~17_combout ))))

	.dataa(\rfile[15][15]~q ),
	.datab(\rfile[14][15]~q ),
	.datac(instruction_D_22),
	.datad(\Mux16~17_combout ),
	.cin(gnd),
	.combout(\Mux16~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~18 .lut_mask = 16'hAFC0;
defparam \Mux16~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N8
cycloneive_lcell_comb \Mux16~10 (
// Equation(s):
// \Mux16~10_combout  = (instruction_D[22] & (((\rfile[10][15]~q ) # (instruction_D[21])))) # (!instruction_D[22] & (\rfile[8][15]~q  & ((!instruction_D[21]))))

	.dataa(\rfile[8][15]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[10][15]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~10 .lut_mask = 16'hCCE2;
defparam \Mux16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N8
cycloneive_lcell_comb \Mux16~11 (
// Equation(s):
// \Mux16~11_combout  = (instruction_D[21] & ((\Mux16~10_combout  & ((\rfile[11][15]~q ))) # (!\Mux16~10_combout  & (\rfile[9][15]~q )))) # (!instruction_D[21] & (((\Mux16~10_combout ))))

	.dataa(\rfile[9][15]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[11][15]~q ),
	.datad(\Mux16~10_combout ),
	.cin(gnd),
	.combout(\Mux16~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~11 .lut_mask = 16'hF388;
defparam \Mux16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N24
cycloneive_lcell_comb \Mux16~14 (
// Equation(s):
// \Mux16~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][15]~q )) # (!instruction_D[22] & ((\rfile[1][15]~q )))))

	.dataa(\rfile[3][15]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[1][15]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux16~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~14 .lut_mask = 16'hB800;
defparam \Mux16~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N10
cycloneive_lcell_comb \Mux16~15 (
// Equation(s):
// \Mux16~15_combout  = (\Mux16~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][15]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux16~14_combout ),
	.datad(\rfile[2][15]~q ),
	.cin(gnd),
	.combout(\Mux16~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~15 .lut_mask = 16'hF2F0;
defparam \Mux16~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N14
cycloneive_lcell_comb \Mux16~12 (
// Equation(s):
// \Mux16~12_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[5][15]~q ))) # (!instruction_D[21] & (\rfile[4][15]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[4][15]~q ),
	.datad(\rfile[5][15]~q ),
	.cin(gnd),
	.combout(\Mux16~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~12 .lut_mask = 16'hDC98;
defparam \Mux16~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N24
cycloneive_lcell_comb \Mux16~13 (
// Equation(s):
// \Mux16~13_combout  = (instruction_D[22] & ((\Mux16~12_combout  & ((\rfile[7][15]~q ))) # (!\Mux16~12_combout  & (\rfile[6][15]~q )))) # (!instruction_D[22] & (((\Mux16~12_combout ))))

	.dataa(\rfile[6][15]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[7][15]~q ),
	.datad(\Mux16~12_combout ),
	.cin(gnd),
	.combout(\Mux16~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~13 .lut_mask = 16'hF388;
defparam \Mux16~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N18
cycloneive_lcell_comb \Mux16~16 (
// Equation(s):
// \Mux16~16_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\Mux16~13_combout )))) # (!instruction_D[23] & (!instruction_D[24] & (\Mux16~15_combout )))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux16~15_combout ),
	.datad(\Mux16~13_combout ),
	.cin(gnd),
	.combout(\Mux16~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~16 .lut_mask = 16'hBA98;
defparam \Mux16~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N14
cycloneive_lcell_comb \Mux17~7 (
// Equation(s):
// \Mux17~7_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[27][14]~q )) # (!instruction_D[24] & ((\rfile[19][14]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[27][14]~q ),
	.datad(\rfile[19][14]~q ),
	.cin(gnd),
	.combout(\Mux17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~7 .lut_mask = 16'hD9C8;
defparam \Mux17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N26
cycloneive_lcell_comb \Mux17~8 (
// Equation(s):
// \Mux17~8_combout  = (instruction_D[23] & ((\Mux17~7_combout  & ((\rfile[31][14]~q ))) # (!\Mux17~7_combout  & (\rfile[23][14]~q )))) # (!instruction_D[23] & (((\Mux17~7_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[23][14]~q ),
	.datac(\rfile[31][14]~q ),
	.datad(\Mux17~7_combout ),
	.cin(gnd),
	.combout(\Mux17~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~8 .lut_mask = 16'hF588;
defparam \Mux17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N18
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[22][14]~q )) # (!instruction_D[23] & ((\rfile[18][14]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[22][14]~q ),
	.datad(\rfile[18][14]~q ),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hD9C8;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N8
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (instruction_D[24] & ((\Mux17~2_combout  & ((\rfile[30][14]~q ))) # (!\Mux17~2_combout  & (\rfile[26][14]~q )))) # (!instruction_D[24] & (((\Mux17~2_combout ))))

	.dataa(\rfile[26][14]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[30][14]~q ),
	.datad(\Mux17~2_combout ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'hF388;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y30_N7
dffeas \rfile[24][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][14] .is_wysiwyg = "true";
defparam \rfile[24][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N20
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (instruction_D[23] & (((\rfile[20][14]~q ) # (instruction_D[24])))) # (!instruction_D[23] & (\rfile[16][14]~q  & ((!instruction_D[24]))))

	.dataa(\rfile[16][14]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[20][14]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hCCE2;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N6
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// \Mux17~5_combout  = (instruction_D[24] & ((\Mux17~4_combout  & (\rfile[28][14]~q )) # (!\Mux17~4_combout  & ((\rfile[24][14]~q ))))) # (!instruction_D[24] & (((\Mux17~4_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[28][14]~q ),
	.datac(\rfile[24][14]~q ),
	.datad(\Mux17~4_combout ),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hDDA0;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N22
cycloneive_lcell_comb \Mux17~6 (
// Equation(s):
// \Mux17~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\Mux17~3_combout )) # (!instruction_D[22] & ((\Mux17~5_combout )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux17~3_combout ),
	.datad(\Mux17~5_combout ),
	.cin(gnd),
	.combout(\Mux17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~6 .lut_mask = 16'hD9C8;
defparam \Mux17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N24
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\rfile[25][14]~q ))) # (!instruction_D[24] & (\rfile[17][14]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[17][14]~q ),
	.datad(\rfile[25][14]~q ),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hDC98;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N10
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (instruction_D[23] & ((\Mux17~0_combout  & ((\rfile[29][14]~q ))) # (!\Mux17~0_combout  & (\rfile[21][14]~q )))) # (!instruction_D[23] & (((\Mux17~0_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[21][14]~q ),
	.datac(\Mux17~0_combout ),
	.datad(\rfile[29][14]~q ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hF858;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N20
cycloneive_lcell_comb \Mux17~10 (
// Equation(s):
// \Mux17~10_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[5][14]~q ))) # (!instruction_D[21] & (\rfile[4][14]~q ))))

	.dataa(instruction_D_22),
	.datab(\rfile[4][14]~q ),
	.datac(instruction_D_21),
	.datad(\rfile[5][14]~q ),
	.cin(gnd),
	.combout(\Mux17~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~10 .lut_mask = 16'hF4A4;
defparam \Mux17~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N26
cycloneive_lcell_comb \Mux17~11 (
// Equation(s):
// \Mux17~11_combout  = (instruction_D[22] & ((\Mux17~10_combout  & (\rfile[7][14]~q )) # (!\Mux17~10_combout  & ((\rfile[6][14]~q ))))) # (!instruction_D[22] & (\Mux17~10_combout ))

	.dataa(instruction_D_22),
	.datab(\Mux17~10_combout ),
	.datac(\rfile[7][14]~q ),
	.datad(\rfile[6][14]~q ),
	.cin(gnd),
	.combout(\Mux17~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~11 .lut_mask = 16'hE6C4;
defparam \Mux17~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N12
cycloneive_lcell_comb \Mux17~17 (
// Equation(s):
// \Mux17~17_combout  = (instruction_D[21] & (((instruction_D[22]) # (\rfile[13][14]~q )))) # (!instruction_D[21] & (\rfile[12][14]~q  & (!instruction_D[22])))

	.dataa(\rfile[12][14]~q ),
	.datab(instruction_D_21),
	.datac(instruction_D_22),
	.datad(\rfile[13][14]~q ),
	.cin(gnd),
	.combout(\Mux17~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~17 .lut_mask = 16'hCEC2;
defparam \Mux17~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N22
cycloneive_lcell_comb \Mux17~18 (
// Equation(s):
// \Mux17~18_combout  = (instruction_D[22] & ((\Mux17~17_combout  & (\rfile[15][14]~q )) # (!\Mux17~17_combout  & ((\rfile[14][14]~q ))))) # (!instruction_D[22] & (((\Mux17~17_combout ))))

	.dataa(\rfile[15][14]~q ),
	.datab(\rfile[14][14]~q ),
	.datac(instruction_D_22),
	.datad(\Mux17~17_combout ),
	.cin(gnd),
	.combout(\Mux17~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~18 .lut_mask = 16'hAFC0;
defparam \Mux17~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N2
cycloneive_lcell_comb \Mux17~14 (
// Equation(s):
// \Mux17~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][14]~q )) # (!instruction_D[22] & ((\rfile[1][14]~q )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[3][14]~q ),
	.datad(\rfile[1][14]~q ),
	.cin(gnd),
	.combout(\Mux17~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~14 .lut_mask = 16'hA280;
defparam \Mux17~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N8
cycloneive_lcell_comb \Mux17~15 (
// Equation(s):
// \Mux17~15_combout  = (\Mux17~14_combout ) # ((!instruction_D[21] & (\rfile[2][14]~q  & instruction_D[22])))

	.dataa(instruction_D_21),
	.datab(\rfile[2][14]~q ),
	.datac(instruction_D_22),
	.datad(\Mux17~14_combout ),
	.cin(gnd),
	.combout(\Mux17~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~15 .lut_mask = 16'hFF40;
defparam \Mux17~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N10
cycloneive_lcell_comb \Mux17~12 (
// Equation(s):
// \Mux17~12_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & ((\rfile[10][14]~q ))) # (!instruction_D[22] & (\rfile[8][14]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[8][14]~q ),
	.datad(\rfile[10][14]~q ),
	.cin(gnd),
	.combout(\Mux17~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~12 .lut_mask = 16'hDC98;
defparam \Mux17~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N4
cycloneive_lcell_comb \Mux17~13 (
// Equation(s):
// \Mux17~13_combout  = (instruction_D[21] & ((\Mux17~12_combout  & (\rfile[11][14]~q )) # (!\Mux17~12_combout  & ((\rfile[9][14]~q ))))) # (!instruction_D[21] & (((\Mux17~12_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[11][14]~q ),
	.datac(\Mux17~12_combout ),
	.datad(\rfile[9][14]~q ),
	.cin(gnd),
	.combout(\Mux17~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~13 .lut_mask = 16'hDAD0;
defparam \Mux17~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N18
cycloneive_lcell_comb \Mux17~16 (
// Equation(s):
// \Mux17~16_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\Mux17~13_combout ))) # (!instruction_D[24] & (\Mux17~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux17~15_combout ),
	.datad(\Mux17~13_combout ),
	.cin(gnd),
	.combout(\Mux17~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~16 .lut_mask = 16'hDC98;
defparam \Mux17~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N10
cycloneive_lcell_comb \Mux18~7 (
// Equation(s):
// \Mux18~7_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[23][13]~q ))) # (!instruction_D[23] & (\rfile[19][13]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[19][13]~q ),
	.datad(\rfile[23][13]~q ),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~7 .lut_mask = 16'hDC98;
defparam \Mux18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y28_N6
cycloneive_lcell_comb \Mux18~8 (
// Equation(s):
// \Mux18~8_combout  = (instruction_D[24] & ((\Mux18~7_combout  & (\rfile[31][13]~q )) # (!\Mux18~7_combout  & ((\rfile[27][13]~q ))))) # (!instruction_D[24] & (((\Mux18~7_combout ))))

	.dataa(\rfile[31][13]~q ),
	.datab(instruction_D_24),
	.datac(\Mux18~7_combout ),
	.datad(\rfile[27][13]~q ),
	.cin(gnd),
	.combout(\Mux18~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~8 .lut_mask = 16'hBCB0;
defparam \Mux18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N24
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[21][13]~q ))) # (!instruction_D[23] & (\rfile[17][13]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[17][13]~q ),
	.datad(\rfile[21][13]~q ),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hDC98;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N26
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (instruction_D[24] & ((\Mux18~0_combout  & ((\rfile[29][13]~q ))) # (!\Mux18~0_combout  & (\rfile[25][13]~q )))) # (!instruction_D[24] & (\Mux18~0_combout ))

	.dataa(instruction_D_24),
	.datab(\Mux18~0_combout ),
	.datac(\rfile[25][13]~q ),
	.datad(\rfile[29][13]~q ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hEC64;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N0
cycloneive_lcell_comb \rfile[20][13]~feeder (
// Equation(s):
// \rfile[20][13]~feeder_combout  = \wdat_WB[13]~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_13),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[20][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[20][13]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[20][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N1
dffeas \rfile[20][13] (
	.clk(!CLK),
	.d(\rfile[20][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][13] .is_wysiwyg = "true";
defparam \rfile[20][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N4
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[24][13]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[16][13]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[16][13]~q ),
	.datad(\rfile[24][13]~q ),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hBA98;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N22
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// \Mux18~5_combout  = (instruction_D[23] & ((\Mux18~4_combout  & ((\rfile[28][13]~q ))) # (!\Mux18~4_combout  & (\rfile[20][13]~q )))) # (!instruction_D[23] & (((\Mux18~4_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[20][13]~q ),
	.datac(\rfile[28][13]~q ),
	.datad(\Mux18~4_combout ),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hF588;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N24
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[26][13]~q )) # (!instruction_D[24] & ((\rfile[18][13]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[26][13]~q ),
	.datad(\rfile[18][13]~q ),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'hD9C8;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N20
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = (instruction_D[23] & ((\Mux18~2_combout  & ((\rfile[30][13]~q ))) # (!\Mux18~2_combout  & (\rfile[22][13]~q )))) # (!instruction_D[23] & (((\Mux18~2_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[22][13]~q ),
	.datac(\rfile[30][13]~q ),
	.datad(\Mux18~2_combout ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'hF588;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N24
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & ((\Mux18~3_combout ))) # (!instruction_D[22] & (\Mux18~5_combout ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux18~5_combout ),
	.datad(\Mux18~3_combout ),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hDC98;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N8
cycloneive_lcell_comb \Mux18~17 (
// Equation(s):
// \Mux18~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][13]~q ))) # (!instruction_D[21] & (\rfile[12][13]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][13]~q ),
	.datad(\rfile[13][13]~q ),
	.cin(gnd),
	.combout(\Mux18~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~17 .lut_mask = 16'hDC98;
defparam \Mux18~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N12
cycloneive_lcell_comb \Mux18~18 (
// Equation(s):
// \Mux18~18_combout  = (instruction_D[22] & ((\Mux18~17_combout  & (\rfile[15][13]~q )) # (!\Mux18~17_combout  & ((\rfile[14][13]~q ))))) # (!instruction_D[22] & (((\Mux18~17_combout ))))

	.dataa(\rfile[15][13]~q ),
	.datab(instruction_D_22),
	.datac(\Mux18~17_combout ),
	.datad(\rfile[14][13]~q ),
	.cin(gnd),
	.combout(\Mux18~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~18 .lut_mask = 16'hBCB0;
defparam \Mux18~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N4
cycloneive_lcell_comb \Mux18~14 (
// Equation(s):
// \Mux18~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][13]~q ))) # (!instruction_D[22] & (\rfile[1][13]~q ))))

	.dataa(instruction_D_21),
	.datab(\rfile[1][13]~q ),
	.datac(instruction_D_22),
	.datad(\rfile[3][13]~q ),
	.cin(gnd),
	.combout(\Mux18~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~14 .lut_mask = 16'hA808;
defparam \Mux18~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y30_N30
cycloneive_lcell_comb \Mux18~15 (
// Equation(s):
// \Mux18~15_combout  = (\Mux18~14_combout ) # ((!instruction_D[21] & (instruction_D[22] & \rfile[2][13]~q )))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux18~14_combout ),
	.datad(\rfile[2][13]~q ),
	.cin(gnd),
	.combout(\Mux18~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~15 .lut_mask = 16'hF4F0;
defparam \Mux18~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N3
dffeas \rfile[7][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][13] .is_wysiwyg = "true";
defparam \rfile[7][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N24
cycloneive_lcell_comb \Mux18~12 (
// Equation(s):
// \Mux18~12_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[5][13]~q )) # (!instruction_D[21] & ((\rfile[4][13]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[5][13]~q ),
	.datad(\rfile[4][13]~q ),
	.cin(gnd),
	.combout(\Mux18~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~12 .lut_mask = 16'hD9C8;
defparam \Mux18~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N2
cycloneive_lcell_comb \Mux18~13 (
// Equation(s):
// \Mux18~13_combout  = (instruction_D[22] & ((\Mux18~12_combout  & ((\rfile[7][13]~q ))) # (!\Mux18~12_combout  & (\rfile[6][13]~q )))) # (!instruction_D[22] & (((\Mux18~12_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[6][13]~q ),
	.datac(\rfile[7][13]~q ),
	.datad(\Mux18~12_combout ),
	.cin(gnd),
	.combout(\Mux18~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~13 .lut_mask = 16'hF588;
defparam \Mux18~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N18
cycloneive_lcell_comb \Mux18~16 (
// Equation(s):
// \Mux18~16_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\Mux18~13_combout ))) # (!instruction_D[23] & (\Mux18~15_combout ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux18~15_combout ),
	.datad(\Mux18~13_combout ),
	.cin(gnd),
	.combout(\Mux18~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~16 .lut_mask = 16'hDC98;
defparam \Mux18~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N20
cycloneive_lcell_comb \Mux18~10 (
// Equation(s):
// \Mux18~10_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\rfile[10][13]~q )) # (!instruction_D[22] & ((\rfile[8][13]~q )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[10][13]~q ),
	.datad(\rfile[8][13]~q ),
	.cin(gnd),
	.combout(\Mux18~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~10 .lut_mask = 16'hD9C8;
defparam \Mux18~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N10
cycloneive_lcell_comb \Mux18~11 (
// Equation(s):
// \Mux18~11_combout  = (instruction_D[21] & ((\Mux18~10_combout  & ((\rfile[11][13]~q ))) # (!\Mux18~10_combout  & (\rfile[9][13]~q )))) # (!instruction_D[21] & (((\Mux18~10_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[9][13]~q ),
	.datac(\rfile[11][13]~q ),
	.datad(\Mux18~10_combout ),
	.cin(gnd),
	.combout(\Mux18~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~11 .lut_mask = 16'hF588;
defparam \Mux18~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N4
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// \Mux19~7_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\rfile[27][12]~q ))) # (!instruction_D[24] & (\rfile[19][12]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[19][12]~q ),
	.datad(\rfile[27][12]~q ),
	.cin(gnd),
	.combout(\Mux19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hDC98;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y29_N30
cycloneive_lcell_comb \Mux19~8 (
// Equation(s):
// \Mux19~8_combout  = (instruction_D[23] & ((\Mux19~7_combout  & (\rfile[31][12]~q )) # (!\Mux19~7_combout  & ((\rfile[23][12]~q ))))) # (!instruction_D[23] & (\Mux19~7_combout ))

	.dataa(instruction_D_23),
	.datab(\Mux19~7_combout ),
	.datac(\rfile[31][12]~q ),
	.datad(\rfile[23][12]~q ),
	.cin(gnd),
	.combout(\Mux19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~8 .lut_mask = 16'hE6C4;
defparam \Mux19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N20
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[25][12]~q )) # (!instruction_D[24] & ((\rfile[17][12]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[25][12]~q ),
	.datad(\rfile[17][12]~q ),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hD9C8;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N24
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (instruction_D[23] & ((\Mux19~0_combout  & (\rfile[29][12]~q )) # (!\Mux19~0_combout  & ((\rfile[21][12]~q ))))) # (!instruction_D[23] & (((\Mux19~0_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[29][12]~q ),
	.datac(\rfile[21][12]~q ),
	.datad(\Mux19~0_combout ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hDDA0;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y36_N23
dffeas \rfile[30][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][12] .is_wysiwyg = "true";
defparam \rfile[30][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N0
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[22][12]~q ))) # (!instruction_D[23] & (\rfile[18][12]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][12]~q ),
	.datad(\rfile[22][12]~q ),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hDC98;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N22
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (instruction_D[24] & ((\Mux19~2_combout  & ((\rfile[30][12]~q ))) # (!\Mux19~2_combout  & (\rfile[26][12]~q )))) # (!instruction_D[24] & (((\Mux19~2_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[26][12]~q ),
	.datac(\rfile[30][12]~q ),
	.datad(\Mux19~2_combout ),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hF588;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y30_N10
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[20][12]~q )))) # (!instruction_D[23] & (!instruction_D[24] & ((\rfile[16][12]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[20][12]~q ),
	.datad(\rfile[16][12]~q ),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'hB9A8;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y30_N23
dffeas \rfile[24][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][12] .is_wysiwyg = "true";
defparam \rfile[24][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N22
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// \Mux19~5_combout  = (instruction_D[24] & ((\Mux19~4_combout  & ((\rfile[28][12]~q ))) # (!\Mux19~4_combout  & (\rfile[24][12]~q )))) # (!instruction_D[24] & (\Mux19~4_combout ))

	.dataa(instruction_D_24),
	.datab(\Mux19~4_combout ),
	.datac(\rfile[24][12]~q ),
	.datad(\rfile[28][12]~q ),
	.cin(gnd),
	.combout(\Mux19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hEC64;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N6
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// \Mux19~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\Mux19~3_combout )) # (!instruction_D[22] & ((\Mux19~5_combout )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux19~3_combout ),
	.datad(\Mux19~5_combout ),
	.cin(gnd),
	.combout(\Mux19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'hD9C8;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N11
dffeas \rfile[4][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][12] .is_wysiwyg = "true";
defparam \rfile[4][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N10
cycloneive_lcell_comb \Mux19~10 (
// Equation(s):
// \Mux19~10_combout  = (instruction_D[21] & ((\rfile[5][12]~q ) # ((instruction_D[22])))) # (!instruction_D[21] & (((\rfile[4][12]~q  & !instruction_D[22]))))

	.dataa(instruction_D_21),
	.datab(\rfile[5][12]~q ),
	.datac(\rfile[4][12]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux19~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~10 .lut_mask = 16'hAAD8;
defparam \Mux19~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N20
cycloneive_lcell_comb \Mux19~11 (
// Equation(s):
// \Mux19~11_combout  = (\Mux19~10_combout  & (((\rfile[7][12]~q ) # (!instruction_D[22])))) # (!\Mux19~10_combout  & (\rfile[6][12]~q  & ((instruction_D[22]))))

	.dataa(\rfile[6][12]~q ),
	.datab(\Mux19~10_combout ),
	.datac(\rfile[7][12]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux19~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~11 .lut_mask = 16'hE2CC;
defparam \Mux19~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N2
cycloneive_lcell_comb \Mux19~14 (
// Equation(s):
// \Mux19~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][12]~q ))) # (!instruction_D[22] & (\rfile[1][12]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][12]~q ),
	.datad(\rfile[3][12]~q ),
	.cin(gnd),
	.combout(\Mux19~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~14 .lut_mask = 16'hC840;
defparam \Mux19~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N30
cycloneive_lcell_comb \Mux19~15 (
// Equation(s):
// \Mux19~15_combout  = (\Mux19~14_combout ) # ((!instruction_D[21] & (instruction_D[22] & \rfile[2][12]~q )))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[2][12]~q ),
	.datad(\Mux19~14_combout ),
	.cin(gnd),
	.combout(\Mux19~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~15 .lut_mask = 16'hFF40;
defparam \Mux19~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N5
dffeas \rfile[10][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][12] .is_wysiwyg = "true";
defparam \rfile[10][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N15
dffeas \rfile[8][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][12] .is_wysiwyg = "true";
defparam \rfile[8][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N14
cycloneive_lcell_comb \Mux19~12 (
// Equation(s):
// \Mux19~12_combout  = (instruction_D[21] & (((instruction_D[22])))) # (!instruction_D[21] & ((instruction_D[22] & (\rfile[10][12]~q )) # (!instruction_D[22] & ((\rfile[8][12]~q )))))

	.dataa(instruction_D_21),
	.datab(\rfile[10][12]~q ),
	.datac(\rfile[8][12]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux19~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~12 .lut_mask = 16'hEE50;
defparam \Mux19~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N18
cycloneive_lcell_comb \Mux19~13 (
// Equation(s):
// \Mux19~13_combout  = (instruction_D[21] & ((\Mux19~12_combout  & ((\rfile[11][12]~q ))) # (!\Mux19~12_combout  & (\rfile[9][12]~q )))) # (!instruction_D[21] & (((\Mux19~12_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[9][12]~q ),
	.datac(\rfile[11][12]~q ),
	.datad(\Mux19~12_combout ),
	.cin(gnd),
	.combout(\Mux19~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~13 .lut_mask = 16'hF588;
defparam \Mux19~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N4
cycloneive_lcell_comb \Mux19~16 (
// Equation(s):
// \Mux19~16_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\Mux19~13_combout ))) # (!instruction_D[24] & (\Mux19~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux19~15_combout ),
	.datad(\Mux19~13_combout ),
	.cin(gnd),
	.combout(\Mux19~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~16 .lut_mask = 16'hDC98;
defparam \Mux19~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N22
cycloneive_lcell_comb \Mux19~17 (
// Equation(s):
// \Mux19~17_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][12]~q )) # (!instruction_D[21] & ((\rfile[12][12]~q )))))

	.dataa(\rfile[13][12]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[12][12]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux19~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~17 .lut_mask = 16'hEE30;
defparam \Mux19~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N28
cycloneive_lcell_comb \Mux19~18 (
// Equation(s):
// \Mux19~18_combout  = (instruction_D[22] & ((\Mux19~17_combout  & (\rfile[15][12]~q )) # (!\Mux19~17_combout  & ((\rfile[14][12]~q ))))) # (!instruction_D[22] & (((\Mux19~17_combout ))))

	.dataa(\rfile[15][12]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[14][12]~q ),
	.datad(\Mux19~17_combout ),
	.cin(gnd),
	.combout(\Mux19~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~18 .lut_mask = 16'hBBC0;
defparam \Mux19~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N0
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[21][11]~q )) # (!instruction_D[23] & ((\rfile[17][11]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[21][11]~q ),
	.datad(\rfile[17][11]~q ),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hD9C8;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y29_N26
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (instruction_D[24] & ((\Mux20~0_combout  & ((\rfile[29][11]~q ))) # (!\Mux20~0_combout  & (\rfile[25][11]~q )))) # (!instruction_D[24] & (((\Mux20~0_combout ))))

	.dataa(\rfile[25][11]~q ),
	.datab(\rfile[29][11]~q ),
	.datac(instruction_D_24),
	.datad(\Mux20~0_combout ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hCFA0;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N10
cycloneive_lcell_comb \Mux20~7 (
// Equation(s):
// \Mux20~7_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[23][11]~q )))) # (!instruction_D[23] & (!instruction_D[24] & ((\rfile[19][11]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[23][11]~q ),
	.datad(\rfile[19][11]~q ),
	.cin(gnd),
	.combout(\Mux20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~7 .lut_mask = 16'hB9A8;
defparam \Mux20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N6
cycloneive_lcell_comb \Mux20~8 (
// Equation(s):
// \Mux20~8_combout  = (instruction_D[24] & ((\Mux20~7_combout  & ((\rfile[31][11]~q ))) # (!\Mux20~7_combout  & (\rfile[27][11]~q )))) # (!instruction_D[24] & (((\Mux20~7_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[27][11]~q ),
	.datac(\rfile[31][11]~q ),
	.datad(\Mux20~7_combout ),
	.cin(gnd),
	.combout(\Mux20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~8 .lut_mask = 16'hF588;
defparam \Mux20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N14
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[24][11]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[16][11]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[24][11]~q ),
	.datad(\rfile[16][11]~q ),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hB9A8;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N24
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// \Mux20~5_combout  = (instruction_D[23] & ((\Mux20~4_combout  & ((\rfile[28][11]~q ))) # (!\Mux20~4_combout  & (\rfile[20][11]~q )))) # (!instruction_D[23] & (((\Mux20~4_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[20][11]~q ),
	.datac(\rfile[28][11]~q ),
	.datad(\Mux20~4_combout ),
	.cin(gnd),
	.combout(\Mux20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hF588;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N26
cycloneive_lcell_comb \rfile[26][11]~feeder (
// Equation(s):
// \rfile[26][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[26][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[26][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[26][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y36_N27
dffeas \rfile[26][11] (
	.clk(!CLK),
	.d(\rfile[26][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][11] .is_wysiwyg = "true";
defparam \rfile[26][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N4
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][11]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[18][11]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][11]~q ),
	.datad(\rfile[26][11]~q ),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hBA98;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N26
cycloneive_lcell_comb \rfile[30][11]~feeder (
// Equation(s):
// \rfile[30][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_11),
	.cin(gnd),
	.combout(\rfile[30][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[30][11]~feeder .lut_mask = 16'hFF00;
defparam \rfile[30][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N27
dffeas \rfile[30][11] (
	.clk(!CLK),
	.d(\rfile[30][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][11] .is_wysiwyg = "true";
defparam \rfile[30][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N22
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (instruction_D[23] & ((\Mux20~2_combout  & ((\rfile[30][11]~q ))) # (!\Mux20~2_combout  & (\rfile[22][11]~q )))) # (!instruction_D[23] & (((\Mux20~2_combout ))))

	.dataa(\rfile[22][11]~q ),
	.datab(instruction_D_23),
	.datac(\Mux20~2_combout ),
	.datad(\rfile[30][11]~q ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'hF838;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N16
cycloneive_lcell_comb \Mux20~6 (
// Equation(s):
// \Mux20~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux20~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & (\Mux20~5_combout )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux20~5_combout ),
	.datad(\Mux20~3_combout ),
	.cin(gnd),
	.combout(\Mux20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~6 .lut_mask = 16'hBA98;
defparam \Mux20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N20
cycloneive_lcell_comb \Mux20~17 (
// Equation(s):
// \Mux20~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][11]~q )) # (!instruction_D[21] & ((\rfile[12][11]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[13][11]~q ),
	.datad(\rfile[12][11]~q ),
	.cin(gnd),
	.combout(\Mux20~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~17 .lut_mask = 16'hD9C8;
defparam \Mux20~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N26
cycloneive_lcell_comb \Mux20~18 (
// Equation(s):
// \Mux20~18_combout  = (instruction_D[22] & ((\Mux20~17_combout  & (\rfile[15][11]~q )) # (!\Mux20~17_combout  & ((\rfile[14][11]~q ))))) # (!instruction_D[22] & (((\Mux20~17_combout ))))

	.dataa(\rfile[15][11]~q ),
	.datab(\rfile[14][11]~q ),
	.datac(instruction_D_22),
	.datad(\Mux20~17_combout ),
	.cin(gnd),
	.combout(\Mux20~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~18 .lut_mask = 16'hAFC0;
defparam \Mux20~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N14
cycloneive_lcell_comb \Mux20~12 (
// Equation(s):
// \Mux20~12_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[5][11]~q ))) # (!instruction_D[21] & (\rfile[4][11]~q ))))

	.dataa(instruction_D_22),
	.datab(\rfile[4][11]~q ),
	.datac(\rfile[5][11]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux20~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~12 .lut_mask = 16'hFA44;
defparam \Mux20~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N12
cycloneive_lcell_comb \rfile[6][11]~feeder (
// Equation(s):
// \rfile[6][11]~feeder_combout  = \wdat_WB[11]~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_11),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[6][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][11]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[6][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N13
dffeas \rfile[6][11] (
	.clk(!CLK),
	.d(\rfile[6][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][11] .is_wysiwyg = "true";
defparam \rfile[6][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N30
cycloneive_lcell_comb \Mux20~13 (
// Equation(s):
// \Mux20~13_combout  = (instruction_D[22] & ((\Mux20~12_combout  & (\rfile[7][11]~q )) # (!\Mux20~12_combout  & ((\rfile[6][11]~q ))))) # (!instruction_D[22] & (((\Mux20~12_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[7][11]~q ),
	.datac(\Mux20~12_combout ),
	.datad(\rfile[6][11]~q ),
	.cin(gnd),
	.combout(\Mux20~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~13 .lut_mask = 16'hDAD0;
defparam \Mux20~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N20
cycloneive_lcell_comb \Mux20~14 (
// Equation(s):
// \Mux20~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][11]~q ))) # (!instruction_D[22] & (\rfile[1][11]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][11]~q ),
	.datad(\rfile[3][11]~q ),
	.cin(gnd),
	.combout(\Mux20~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~14 .lut_mask = 16'hC840;
defparam \Mux20~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N14
cycloneive_lcell_comb \Mux20~15 (
// Equation(s):
// \Mux20~15_combout  = (\Mux20~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][11]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[2][11]~q ),
	.datad(\Mux20~14_combout ),
	.cin(gnd),
	.combout(\Mux20~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~15 .lut_mask = 16'hFF20;
defparam \Mux20~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N8
cycloneive_lcell_comb \Mux20~16 (
// Equation(s):
// \Mux20~16_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\Mux20~13_combout )) # (!instruction_D[23] & ((\Mux20~15_combout )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux20~13_combout ),
	.datad(\Mux20~15_combout ),
	.cin(gnd),
	.combout(\Mux20~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~16 .lut_mask = 16'hD9C8;
defparam \Mux20~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N6
cycloneive_lcell_comb \Mux20~10 (
// Equation(s):
// \Mux20~10_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & ((\rfile[10][11]~q ))) # (!instruction_D[22] & (\rfile[8][11]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[8][11]~q ),
	.datad(\rfile[10][11]~q ),
	.cin(gnd),
	.combout(\Mux20~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~10 .lut_mask = 16'hDC98;
defparam \Mux20~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N28
cycloneive_lcell_comb \Mux20~11 (
// Equation(s):
// \Mux20~11_combout  = (\Mux20~10_combout  & (((\rfile[11][11]~q )) # (!instruction_D[21]))) # (!\Mux20~10_combout  & (instruction_D[21] & ((\rfile[9][11]~q ))))

	.dataa(\Mux20~10_combout ),
	.datab(instruction_D_21),
	.datac(\rfile[11][11]~q ),
	.datad(\rfile[9][11]~q ),
	.cin(gnd),
	.combout(\Mux20~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~11 .lut_mask = 16'hE6A2;
defparam \Mux20~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N31
dffeas \rfile[17][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][10] .is_wysiwyg = "true";
defparam \rfile[17][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N30
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[25][10]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[17][10]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[17][10]~q ),
	.datad(\rfile[25][10]~q ),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hBA98;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N8
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (\Mux21~0_combout  & (((\rfile[29][10]~q )) # (!instruction_D[23]))) # (!\Mux21~0_combout  & (instruction_D[23] & (\rfile[21][10]~q )))

	.dataa(\Mux21~0_combout ),
	.datab(instruction_D_23),
	.datac(\rfile[21][10]~q ),
	.datad(\rfile[29][10]~q ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hEA62;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N24
cycloneive_lcell_comb \Mux21~7 (
// Equation(s):
// \Mux21~7_combout  = (instruction_D[24] & (((instruction_D[23]) # (\rfile[27][10]~q )))) # (!instruction_D[24] & (\rfile[19][10]~q  & (!instruction_D[23])))

	.dataa(instruction_D_24),
	.datab(\rfile[19][10]~q ),
	.datac(instruction_D_23),
	.datad(\rfile[27][10]~q ),
	.cin(gnd),
	.combout(\Mux21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~7 .lut_mask = 16'hAEA4;
defparam \Mux21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N22
cycloneive_lcell_comb \Mux21~8 (
// Equation(s):
// \Mux21~8_combout  = (instruction_D[23] & ((\Mux21~7_combout  & ((\rfile[31][10]~q ))) # (!\Mux21~7_combout  & (\rfile[23][10]~q )))) # (!instruction_D[23] & (((\Mux21~7_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[23][10]~q ),
	.datac(\rfile[31][10]~q ),
	.datad(\Mux21~7_combout ),
	.cin(gnd),
	.combout(\Mux21~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~8 .lut_mask = 16'hF588;
defparam \Mux21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N4
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// \Mux21~5_combout  = (\Mux21~4_combout  & (((\rfile[28][10]~q ) # (!instruction_D[24])))) # (!\Mux21~4_combout  & (\rfile[24][10]~q  & ((instruction_D[24]))))

	.dataa(\Mux21~4_combout ),
	.datab(\rfile[24][10]~q ),
	.datac(\rfile[28][10]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hE4AA;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y36_N11
dffeas \rfile[26][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][10] .is_wysiwyg = "true";
defparam \rfile[26][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y36_N4
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[22][10]~q )))) # (!instruction_D[23] & (!instruction_D[24] & (\rfile[18][10]~q )))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[18][10]~q ),
	.datad(\rfile[22][10]~q ),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hBA98;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N10
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (instruction_D[24] & ((\Mux21~2_combout  & (\rfile[30][10]~q )) # (!\Mux21~2_combout  & ((\rfile[26][10]~q ))))) # (!instruction_D[24] & (((\Mux21~2_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[30][10]~q ),
	.datac(\rfile[26][10]~q ),
	.datad(\Mux21~2_combout ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'hDDA0;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N6
cycloneive_lcell_comb \Mux21~6 (
// Equation(s):
// \Mux21~6_combout  = (instruction_D[22] & (((instruction_D[21]) # (\Mux21~3_combout )))) # (!instruction_D[22] & (\Mux21~5_combout  & (!instruction_D[21])))

	.dataa(\Mux21~5_combout ),
	.datab(instruction_D_22),
	.datac(instruction_D_21),
	.datad(\Mux21~3_combout ),
	.cin(gnd),
	.combout(\Mux21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~6 .lut_mask = 16'hCEC2;
defparam \Mux21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N8
cycloneive_lcell_comb \Mux21~10 (
// Equation(s):
// \Mux21~10_combout  = (instruction_D[21] & ((instruction_D[22]) # ((\rfile[5][10]~q )))) # (!instruction_D[21] & (!instruction_D[22] & ((\rfile[4][10]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[5][10]~q ),
	.datad(\rfile[4][10]~q ),
	.cin(gnd),
	.combout(\Mux21~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~10 .lut_mask = 16'hB9A8;
defparam \Mux21~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N20
cycloneive_lcell_comb \Mux21~11 (
// Equation(s):
// \Mux21~11_combout  = (\Mux21~10_combout  & (((\rfile[7][10]~q )) # (!instruction_D[22]))) # (!\Mux21~10_combout  & (instruction_D[22] & (\rfile[6][10]~q )))

	.dataa(\Mux21~10_combout ),
	.datab(instruction_D_22),
	.datac(\rfile[6][10]~q ),
	.datad(\rfile[7][10]~q ),
	.cin(gnd),
	.combout(\Mux21~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~11 .lut_mask = 16'hEA62;
defparam \Mux21~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N18
cycloneive_lcell_comb \Mux21~17 (
// Equation(s):
// \Mux21~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][10]~q ))) # (!instruction_D[21] & (\rfile[12][10]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][10]~q ),
	.datad(\rfile[13][10]~q ),
	.cin(gnd),
	.combout(\Mux21~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~17 .lut_mask = 16'hDC98;
defparam \Mux21~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N14
cycloneive_lcell_comb \Mux21~18 (
// Equation(s):
// \Mux21~18_combout  = (instruction_D[22] & ((\Mux21~17_combout  & (\rfile[15][10]~q )) # (!\Mux21~17_combout  & ((\rfile[14][10]~q ))))) # (!instruction_D[22] & (((\Mux21~17_combout ))))

	.dataa(\rfile[15][10]~q ),
	.datab(\rfile[14][10]~q ),
	.datac(instruction_D_22),
	.datad(\Mux21~17_combout ),
	.cin(gnd),
	.combout(\Mux21~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~18 .lut_mask = 16'hAFC0;
defparam \Mux21~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N22
cycloneive_lcell_comb \Mux21~13 (
// Equation(s):
// \Mux21~13_combout  = (\Mux21~12_combout  & ((\rfile[11][10]~q ) # ((!instruction_D[21])))) # (!\Mux21~12_combout  & (((\rfile[9][10]~q  & instruction_D[21]))))

	.dataa(\Mux21~12_combout ),
	.datab(\rfile[11][10]~q ),
	.datac(\rfile[9][10]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux21~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~13 .lut_mask = 16'hD8AA;
defparam \Mux21~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N26
cycloneive_lcell_comb \Mux21~14 (
// Equation(s):
// \Mux21~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][10]~q )) # (!instruction_D[22] & ((\rfile[1][10]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[3][10]~q ),
	.datad(\rfile[1][10]~q ),
	.cin(gnd),
	.combout(\Mux21~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~14 .lut_mask = 16'hC480;
defparam \Mux21~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N20
cycloneive_lcell_comb \Mux21~15 (
// Equation(s):
// \Mux21~15_combout  = (\Mux21~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][10]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[2][10]~q ),
	.datad(\Mux21~14_combout ),
	.cin(gnd),
	.combout(\Mux21~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~15 .lut_mask = 16'hFF20;
defparam \Mux21~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N30
cycloneive_lcell_comb \Mux21~16 (
// Equation(s):
// \Mux21~16_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\Mux21~13_combout )))) # (!instruction_D[24] & (!instruction_D[23] & ((\Mux21~15_combout ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux21~13_combout ),
	.datad(\Mux21~15_combout ),
	.cin(gnd),
	.combout(\Mux21~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~16 .lut_mask = 16'hB9A8;
defparam \Mux21~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y32_N13
dffeas \rfile[20][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][9] .is_wysiwyg = "true";
defparam \rfile[20][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N6
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[24][9]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[16][9]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[24][9]~q ),
	.datad(\rfile[16][9]~q ),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hB9A8;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N12
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// \Mux22~5_combout  = (instruction_D[23] & ((\Mux22~4_combout  & (\rfile[28][9]~q )) # (!\Mux22~4_combout  & ((\rfile[20][9]~q ))))) # (!instruction_D[23] & (((\Mux22~4_combout ))))

	.dataa(\rfile[28][9]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[20][9]~q ),
	.datad(\Mux22~4_combout ),
	.cin(gnd),
	.combout(\Mux22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hBBC0;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N28
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][9]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[18][9]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][9]~q ),
	.datad(\rfile[26][9]~q ),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hBA98;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N10
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (\Mux22~2_combout  & (((\rfile[30][9]~q ) # (!instruction_D[23])))) # (!\Mux22~2_combout  & (\rfile[22][9]~q  & ((instruction_D[23]))))

	.dataa(\rfile[22][9]~q ),
	.datab(\rfile[30][9]~q ),
	.datac(\Mux22~2_combout ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'hCAF0;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N12
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// \Mux22~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & ((\Mux22~3_combout ))) # (!instruction_D[22] & (\Mux22~5_combout ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux22~5_combout ),
	.datad(\Mux22~3_combout ),
	.cin(gnd),
	.combout(\Mux22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'hDC98;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N10
cycloneive_lcell_comb \Mux22~7 (
// Equation(s):
// \Mux22~7_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[23][9]~q ))) # (!instruction_D[23] & (\rfile[19][9]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[19][9]~q ),
	.datad(\rfile[23][9]~q ),
	.cin(gnd),
	.combout(\Mux22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~7 .lut_mask = 16'hDC98;
defparam \Mux22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N26
cycloneive_lcell_comb \Mux22~8 (
// Equation(s):
// \Mux22~8_combout  = (instruction_D[24] & ((\Mux22~7_combout  & ((\rfile[31][9]~q ))) # (!\Mux22~7_combout  & (\rfile[27][9]~q )))) # (!instruction_D[24] & (((\Mux22~7_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[27][9]~q ),
	.datac(\rfile[31][9]~q ),
	.datad(\Mux22~7_combout ),
	.cin(gnd),
	.combout(\Mux22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~8 .lut_mask = 16'hF588;
defparam \Mux22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N4
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[21][9]~q )) # (!instruction_D[23] & ((\rfile[17][9]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[21][9]~q ),
	.datad(\rfile[17][9]~q ),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hD9C8;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N6
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (instruction_D[24] & ((\Mux22~0_combout  & (\rfile[29][9]~q )) # (!\Mux22~0_combout  & ((\rfile[25][9]~q ))))) # (!instruction_D[24] & (((\Mux22~0_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[29][9]~q ),
	.datac(\rfile[25][9]~q ),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hDDA0;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N12
cycloneive_lcell_comb \Mux22~10 (
// Equation(s):
// \Mux22~10_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\rfile[10][9]~q )) # (!instruction_D[22] & ((\rfile[8][9]~q )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[10][9]~q ),
	.datad(\rfile[8][9]~q ),
	.cin(gnd),
	.combout(\Mux22~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~10 .lut_mask = 16'hD9C8;
defparam \Mux22~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N30
cycloneive_lcell_comb \Mux22~11 (
// Equation(s):
// \Mux22~11_combout  = (instruction_D[21] & ((\Mux22~10_combout  & (\rfile[11][9]~q )) # (!\Mux22~10_combout  & ((\rfile[9][9]~q ))))) # (!instruction_D[21] & (\Mux22~10_combout ))

	.dataa(instruction_D_21),
	.datab(\Mux22~10_combout ),
	.datac(\rfile[11][9]~q ),
	.datad(\rfile[9][9]~q ),
	.cin(gnd),
	.combout(\Mux22~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~11 .lut_mask = 16'hE6C4;
defparam \Mux22~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N9
dffeas \rfile[4][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][9] .is_wysiwyg = "true";
defparam \rfile[4][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N27
dffeas \rfile[5][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][9] .is_wysiwyg = "true";
defparam \rfile[5][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N8
cycloneive_lcell_comb \Mux22~12 (
// Equation(s):
// \Mux22~12_combout  = (instruction_D[21] & ((instruction_D[22]) # ((\rfile[5][9]~q )))) # (!instruction_D[21] & (!instruction_D[22] & (\rfile[4][9]~q )))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[4][9]~q ),
	.datad(\rfile[5][9]~q ),
	.cin(gnd),
	.combout(\Mux22~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~12 .lut_mask = 16'hBA98;
defparam \Mux22~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N30
cycloneive_lcell_comb \Mux22~13 (
// Equation(s):
// \Mux22~13_combout  = (\Mux22~12_combout  & (((\rfile[7][9]~q ) # (!instruction_D[22])))) # (!\Mux22~12_combout  & (\rfile[6][9]~q  & ((instruction_D[22]))))

	.dataa(\rfile[6][9]~q ),
	.datab(\Mux22~12_combout ),
	.datac(\rfile[7][9]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux22~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~13 .lut_mask = 16'hE2CC;
defparam \Mux22~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N24
cycloneive_lcell_comb \Mux22~14 (
// Equation(s):
// \Mux22~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][9]~q )) # (!instruction_D[22] & ((\rfile[1][9]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[3][9]~q ),
	.datad(\rfile[1][9]~q ),
	.cin(gnd),
	.combout(\Mux22~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~14 .lut_mask = 16'hC480;
defparam \Mux22~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N24
cycloneive_lcell_comb \Mux22~15 (
// Equation(s):
// \Mux22~15_combout  = (\Mux22~14_combout ) # ((\rfile[2][9]~q  & (!instruction_D[21] & instruction_D[22])))

	.dataa(\rfile[2][9]~q ),
	.datab(instruction_D_21),
	.datac(instruction_D_22),
	.datad(\Mux22~14_combout ),
	.cin(gnd),
	.combout(\Mux22~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~15 .lut_mask = 16'hFF20;
defparam \Mux22~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N6
cycloneive_lcell_comb \Mux22~16 (
// Equation(s):
// \Mux22~16_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\Mux22~13_combout )) # (!instruction_D[23] & ((\Mux22~15_combout )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux22~13_combout ),
	.datad(\Mux22~15_combout ),
	.cin(gnd),
	.combout(\Mux22~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~16 .lut_mask = 16'hD9C8;
defparam \Mux22~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N8
cycloneive_lcell_comb \Mux22~17 (
// Equation(s):
// \Mux22~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][9]~q )) # (!instruction_D[21] & ((\rfile[12][9]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[13][9]~q ),
	.datad(\rfile[12][9]~q ),
	.cin(gnd),
	.combout(\Mux22~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~17 .lut_mask = 16'hD9C8;
defparam \Mux22~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N8
cycloneive_lcell_comb \Mux22~18 (
// Equation(s):
// \Mux22~18_combout  = (instruction_D[22] & ((\Mux22~17_combout  & (\rfile[15][9]~q )) # (!\Mux22~17_combout  & ((\rfile[14][9]~q ))))) # (!instruction_D[22] & (((\Mux22~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[15][9]~q ),
	.datac(\rfile[14][9]~q ),
	.datad(\Mux22~17_combout ),
	.cin(gnd),
	.combout(\Mux22~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~18 .lut_mask = 16'hDDA0;
defparam \Mux22~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N2
cycloneive_lcell_comb \Mux59~7 (
// Equation(s):
// \Mux59~7_combout  = (instruction_D[19] & ((instruction_D[18]) # ((\rfile[27][4]~q )))) # (!instruction_D[19] & (!instruction_D[18] & (\rfile[19][4]~q )))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[19][4]~q ),
	.datad(\rfile[27][4]~q ),
	.cin(gnd),
	.combout(\Mux59~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~7 .lut_mask = 16'hBA98;
defparam \Mux59~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N2
cycloneive_lcell_comb \Mux59~8 (
// Equation(s):
// \Mux59~8_combout  = (instruction_D[18] & ((\Mux59~7_combout  & (\rfile[31][4]~q )) # (!\Mux59~7_combout  & ((\rfile[23][4]~q ))))) # (!instruction_D[18] & (((\Mux59~7_combout ))))

	.dataa(instruction_D_18),
	.datab(\rfile[31][4]~q ),
	.datac(\rfile[23][4]~q ),
	.datad(\Mux59~7_combout ),
	.cin(gnd),
	.combout(\Mux59~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~8 .lut_mask = 16'hDDA0;
defparam \Mux59~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N8
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\rfile[25][4]~q )) # (!instruction_D[19] & ((\rfile[17][4]~q )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\rfile[25][4]~q ),
	.datad(\rfile[17][4]~q ),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'hD9C8;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N12
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (instruction_D[18] & ((\Mux59~0_combout  & ((\rfile[29][4]~q ))) # (!\Mux59~0_combout  & (\rfile[21][4]~q )))) # (!instruction_D[18] & (((\Mux59~0_combout ))))

	.dataa(\rfile[21][4]~q ),
	.datab(instruction_D_18),
	.datac(\rfile[29][4]~q ),
	.datad(\Mux59~0_combout ),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hF388;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y34_N22
cycloneive_lcell_comb \rfile[30][4]~feeder (
// Equation(s):
// \rfile[30][4]~feeder_combout  = \wdat_WB[4]~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_4),
	.cin(gnd),
	.combout(\rfile[30][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[30][4]~feeder .lut_mask = 16'hFF00;
defparam \rfile[30][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y34_N23
dffeas \rfile[30][4] (
	.clk(!CLK),
	.d(\rfile[30][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[30][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[30][4] .is_wysiwyg = "true";
defparam \rfile[30][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N20
cycloneive_lcell_comb \Mux59~2 (
// Equation(s):
// \Mux59~2_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & ((\rfile[22][4]~q ))) # (!instruction_D[18] & (\rfile[18][4]~q ))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[18][4]~q ),
	.datad(\rfile[22][4]~q ),
	.cin(gnd),
	.combout(\Mux59~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~2 .lut_mask = 16'hDC98;
defparam \Mux59~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y34_N30
cycloneive_lcell_comb \Mux59~3 (
// Equation(s):
// \Mux59~3_combout  = (instruction_D[19] & ((\Mux59~2_combout  & ((\rfile[30][4]~q ))) # (!\Mux59~2_combout  & (\rfile[26][4]~q )))) # (!instruction_D[19] & (((\Mux59~2_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[26][4]~q ),
	.datac(\rfile[30][4]~q ),
	.datad(\Mux59~2_combout ),
	.cin(gnd),
	.combout(\Mux59~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~3 .lut_mask = 16'hF588;
defparam \Mux59~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y32_N4
cycloneive_lcell_comb \Mux59~4 (
// Equation(s):
// \Mux59~4_combout  = (instruction_D[19] & (instruction_D[18])) # (!instruction_D[19] & ((instruction_D[18] & (\rfile[20][4]~q )) # (!instruction_D[18] & ((\rfile[16][4]~q )))))

	.dataa(instruction_D_19),
	.datab(instruction_D_18),
	.datac(\rfile[20][4]~q ),
	.datad(\rfile[16][4]~q ),
	.cin(gnd),
	.combout(\Mux59~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~4 .lut_mask = 16'hD9C8;
defparam \Mux59~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N16
cycloneive_lcell_comb \Mux59~5 (
// Equation(s):
// \Mux59~5_combout  = (instruction_D[19] & ((\Mux59~4_combout  & (\rfile[28][4]~q )) # (!\Mux59~4_combout  & ((\rfile[24][4]~q ))))) # (!instruction_D[19] & (((\Mux59~4_combout ))))

	.dataa(instruction_D_19),
	.datab(\rfile[28][4]~q ),
	.datac(\rfile[24][4]~q ),
	.datad(\Mux59~4_combout ),
	.cin(gnd),
	.combout(\Mux59~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~5 .lut_mask = 16'hDDA0;
defparam \Mux59~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N10
cycloneive_lcell_comb \Mux59~6 (
// Equation(s):
// \Mux59~6_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & (\Mux59~3_combout )) # (!instruction_D[17] & ((\Mux59~5_combout )))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\Mux59~3_combout ),
	.datad(\Mux59~5_combout ),
	.cin(gnd),
	.combout(\Mux59~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~6 .lut_mask = 16'hD9C8;
defparam \Mux59~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N2
cycloneive_lcell_comb \Mux59~17 (
// Equation(s):
// \Mux59~17_combout  = (instruction_D[16] & ((instruction_D[17]) # ((\rfile[13][4]~q )))) # (!instruction_D[16] & (!instruction_D[17] & (\rfile[12][4]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[12][4]~q ),
	.datad(\rfile[13][4]~q ),
	.cin(gnd),
	.combout(\Mux59~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~17 .lut_mask = 16'hBA98;
defparam \Mux59~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N0
cycloneive_lcell_comb \Mux59~18 (
// Equation(s):
// \Mux59~18_combout  = (\Mux59~17_combout  & (((\rfile[15][4]~q ) # (!instruction_D[17])))) # (!\Mux59~17_combout  & (\rfile[14][4]~q  & (instruction_D[17])))

	.dataa(\rfile[14][4]~q ),
	.datab(\Mux59~17_combout ),
	.datac(instruction_D_17),
	.datad(\rfile[15][4]~q ),
	.cin(gnd),
	.combout(\Mux59~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~18 .lut_mask = 16'hEC2C;
defparam \Mux59~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N2
cycloneive_lcell_comb \Mux59~12 (
// Equation(s):
// \Mux59~12_combout  = (instruction_D[16] & (instruction_D[17])) # (!instruction_D[16] & ((instruction_D[17] & ((\rfile[10][4]~q ))) # (!instruction_D[17] & (\rfile[8][4]~q ))))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[8][4]~q ),
	.datad(\rfile[10][4]~q ),
	.cin(gnd),
	.combout(\Mux59~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~12 .lut_mask = 16'hDC98;
defparam \Mux59~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N26
cycloneive_lcell_comb \Mux59~13 (
// Equation(s):
// \Mux59~13_combout  = (instruction_D[16] & ((\Mux59~12_combout  & (\rfile[11][4]~q )) # (!\Mux59~12_combout  & ((\rfile[9][4]~q ))))) # (!instruction_D[16] & (((\Mux59~12_combout ))))

	.dataa(instruction_D_16),
	.datab(\rfile[11][4]~q ),
	.datac(\rfile[9][4]~q ),
	.datad(\Mux59~12_combout ),
	.cin(gnd),
	.combout(\Mux59~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~13 .lut_mask = 16'hDDA0;
defparam \Mux59~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N28
cycloneive_lcell_comb \Mux59~14 (
// Equation(s):
// \Mux59~14_combout  = (instruction_D[16] & ((instruction_D[17] & ((\rfile[3][4]~q ))) # (!instruction_D[17] & (\rfile[1][4]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[1][4]~q ),
	.datad(\rfile[3][4]~q ),
	.cin(gnd),
	.combout(\Mux59~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~14 .lut_mask = 16'hC840;
defparam \Mux59~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N28
cycloneive_lcell_comb \Mux59~15 (
// Equation(s):
// \Mux59~15_combout  = (\Mux59~14_combout ) # ((!instruction_D[16] & (instruction_D[17] & \rfile[2][4]~q )))

	.dataa(instruction_D_16),
	.datab(instruction_D_17),
	.datac(\rfile[2][4]~q ),
	.datad(\Mux59~14_combout ),
	.cin(gnd),
	.combout(\Mux59~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~15 .lut_mask = 16'hFF40;
defparam \Mux59~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N22
cycloneive_lcell_comb \Mux59~16 (
// Equation(s):
// \Mux59~16_combout  = (instruction_D[18] & (instruction_D[19])) # (!instruction_D[18] & ((instruction_D[19] & (\Mux59~13_combout )) # (!instruction_D[19] & ((\Mux59~15_combout )))))

	.dataa(instruction_D_18),
	.datab(instruction_D_19),
	.datac(\Mux59~13_combout ),
	.datad(\Mux59~15_combout ),
	.cin(gnd),
	.combout(\Mux59~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~16 .lut_mask = 16'hD9C8;
defparam \Mux59~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N6
cycloneive_lcell_comb \Mux59~10 (
// Equation(s):
// \Mux59~10_combout  = (instruction_D[17] & (instruction_D[16])) # (!instruction_D[17] & ((instruction_D[16] & ((\rfile[5][4]~q ))) # (!instruction_D[16] & (\rfile[4][4]~q ))))

	.dataa(instruction_D_17),
	.datab(instruction_D_16),
	.datac(\rfile[4][4]~q ),
	.datad(\rfile[5][4]~q ),
	.cin(gnd),
	.combout(\Mux59~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~10 .lut_mask = 16'hDC98;
defparam \Mux59~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N14
cycloneive_lcell_comb \Mux59~11 (
// Equation(s):
// \Mux59~11_combout  = (instruction_D[17] & ((\Mux59~10_combout  & ((\rfile[7][4]~q ))) # (!\Mux59~10_combout  & (\rfile[6][4]~q )))) # (!instruction_D[17] & (((\Mux59~10_combout ))))

	.dataa(instruction_D_17),
	.datab(\rfile[6][4]~q ),
	.datac(\rfile[7][4]~q ),
	.datad(\Mux59~10_combout ),
	.cin(gnd),
	.combout(\Mux59~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~11 .lut_mask = 16'hF588;
defparam \Mux59~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N0
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[21][31]~q )))) # (!instruction_D[23] & (!instruction_D[24] & ((\rfile[17][31]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[21][31]~q ),
	.datad(\rfile[17][31]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hB9A8;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N6
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (instruction_D[24] & ((\Mux0~0_combout  & ((\rfile[29][31]~q ))) # (!\Mux0~0_combout  & (\rfile[25][31]~q )))) # (!instruction_D[24] & (((\Mux0~0_combout ))))

	.dataa(\rfile[25][31]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[29][31]~q ),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hF388;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N8
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[24][31]~q )) # (!instruction_D[24] & ((\rfile[16][31]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[24][31]~q ),
	.datad(\rfile[16][31]~q ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'hD9C8;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N1
dffeas \rfile[20][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][31] .is_wysiwyg = "true";
defparam \rfile[20][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N0
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (instruction_D[23] & ((\Mux0~4_combout  & ((\rfile[28][31]~q ))) # (!\Mux0~4_combout  & (\rfile[20][31]~q )))) # (!instruction_D[23] & (\Mux0~4_combout ))

	.dataa(instruction_D_23),
	.datab(\Mux0~4_combout ),
	.datac(\rfile[20][31]~q ),
	.datad(\rfile[28][31]~q ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hEC64;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y36_N17
dffeas \rfile[26][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][31] .is_wysiwyg = "true";
defparam \rfile[26][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y34_N23
dffeas \rfile[18][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][31] .is_wysiwyg = "true";
defparam \rfile[18][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N16
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][31]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[18][31]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[26][31]~q ),
	.datad(\rfile[18][31]~q ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hB9A8;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N14
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (instruction_D[23] & ((\Mux0~2_combout  & ((\rfile[30][31]~q ))) # (!\Mux0~2_combout  & (\rfile[22][31]~q )))) # (!instruction_D[23] & (((\Mux0~2_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[22][31]~q ),
	.datac(\rfile[30][31]~q ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'hF588;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N14
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux0~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & (\Mux0~5_combout )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux0~5_combout ),
	.datad(\Mux0~3_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'hBA98;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N0
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// \Mux0~7_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[23][31]~q )) # (!instruction_D[23] & ((\rfile[19][31]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[23][31]~q ),
	.datad(\rfile[19][31]~q ),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hD9C8;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N4
cycloneive_lcell_comb \Mux0~8 (
// Equation(s):
// \Mux0~8_combout  = (instruction_D[24] & ((\Mux0~7_combout  & (\rfile[31][31]~q )) # (!\Mux0~7_combout  & ((\rfile[27][31]~q ))))) # (!instruction_D[24] & (((\Mux0~7_combout ))))

	.dataa(\rfile[31][31]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[27][31]~q ),
	.datad(\Mux0~7_combout ),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~8 .lut_mask = 16'hBBC0;
defparam \Mux0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N23
dffeas \rfile[8][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[8][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[8][31] .is_wysiwyg = "true";
defparam \rfile[8][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N22
cycloneive_lcell_comb \Mux0~10 (
// Equation(s):
// \Mux0~10_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][31]~q )))) # (!instruction_D[22] & (!instruction_D[21] & (\rfile[8][31]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[8][31]~q ),
	.datad(\rfile[10][31]~q ),
	.cin(gnd),
	.combout(\Mux0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~10 .lut_mask = 16'hBA98;
defparam \Mux0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N2
cycloneive_lcell_comb \Mux0~11 (
// Equation(s):
// \Mux0~11_combout  = (\Mux0~10_combout  & ((\rfile[11][31]~q ) # ((!instruction_D[21])))) # (!\Mux0~10_combout  & (((\rfile[9][31]~q  & instruction_D[21]))))

	.dataa(\rfile[11][31]~q ),
	.datab(\rfile[9][31]~q ),
	.datac(\Mux0~10_combout ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~11 .lut_mask = 16'hACF0;
defparam \Mux0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N4
cycloneive_lcell_comb \Mux0~17 (
// Equation(s):
// \Mux0~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][31]~q )) # (!instruction_D[21] & ((\rfile[12][31]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[13][31]~q ),
	.datad(\rfile[12][31]~q ),
	.cin(gnd),
	.combout(\Mux0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~17 .lut_mask = 16'hD9C8;
defparam \Mux0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N2
cycloneive_lcell_comb \Mux0~18 (
// Equation(s):
// \Mux0~18_combout  = (\Mux0~17_combout  & (((\rfile[15][31]~q )) # (!instruction_D[22]))) # (!\Mux0~17_combout  & (instruction_D[22] & ((\rfile[14][31]~q ))))

	.dataa(\Mux0~17_combout ),
	.datab(instruction_D_22),
	.datac(\rfile[15][31]~q ),
	.datad(\rfile[14][31]~q ),
	.cin(gnd),
	.combout(\Mux0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~18 .lut_mask = 16'hE6A2;
defparam \Mux0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N27
dffeas \rfile[7][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][31] .is_wysiwyg = "true";
defparam \rfile[7][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N27
dffeas \rfile[4][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][31] .is_wysiwyg = "true";
defparam \rfile[4][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N26
cycloneive_lcell_comb \Mux0~12 (
// Equation(s):
// \Mux0~12_combout  = (instruction_D[21] & ((instruction_D[22]) # ((\rfile[5][31]~q )))) # (!instruction_D[21] & (!instruction_D[22] & (\rfile[4][31]~q )))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[4][31]~q ),
	.datad(\rfile[5][31]~q ),
	.cin(gnd),
	.combout(\Mux0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~12 .lut_mask = 16'hBA98;
defparam \Mux0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N26
cycloneive_lcell_comb \Mux0~13 (
// Equation(s):
// \Mux0~13_combout  = (instruction_D[22] & ((\Mux0~12_combout  & ((\rfile[7][31]~q ))) # (!\Mux0~12_combout  & (\rfile[6][31]~q )))) # (!instruction_D[22] & (((\Mux0~12_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[6][31]~q ),
	.datac(\rfile[7][31]~q ),
	.datad(\Mux0~12_combout ),
	.cin(gnd),
	.combout(\Mux0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~13 .lut_mask = 16'hF588;
defparam \Mux0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N28
cycloneive_lcell_comb \Mux0~15 (
// Equation(s):
// \Mux0~15_combout  = (\Mux0~14_combout ) # ((\rfile[2][31]~q  & (!instruction_D[21] & instruction_D[22])))

	.dataa(\Mux0~14_combout ),
	.datab(\rfile[2][31]~q ),
	.datac(instruction_D_21),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~15 .lut_mask = 16'hAEAA;
defparam \Mux0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N6
cycloneive_lcell_comb \Mux0~16 (
// Equation(s):
// \Mux0~16_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\Mux0~13_combout )) # (!instruction_D[23] & ((\Mux0~15_combout )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux0~13_combout ),
	.datad(\Mux0~15_combout ),
	.cin(gnd),
	.combout(\Mux0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~16 .lut_mask = 16'hD9C8;
defparam \Mux0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N6
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (instruction_D[24] & (((instruction_D[23])))) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[23][29]~q )) # (!instruction_D[23] & ((\rfile[19][29]~q )))))

	.dataa(instruction_D_24),
	.datab(\rfile[23][29]~q ),
	.datac(\rfile[19][29]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hEE50;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N26
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (instruction_D[24] & ((\Mux2~7_combout  & ((\rfile[31][29]~q ))) # (!\Mux2~7_combout  & (\rfile[27][29]~q )))) # (!instruction_D[24] & (((\Mux2~7_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[27][29]~q ),
	.datac(\rfile[31][29]~q ),
	.datad(\Mux2~7_combout ),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hF588;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N14
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[21][29]~q ))) # (!instruction_D[23] & (\rfile[17][29]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[17][29]~q ),
	.datad(\rfile[21][29]~q ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hDC98;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N18
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (instruction_D[24] & ((\Mux2~0_combout  & ((\rfile[29][29]~q ))) # (!\Mux2~0_combout  & (\rfile[25][29]~q )))) # (!instruction_D[24] & (((\Mux2~0_combout ))))

	.dataa(\rfile[25][29]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[29][29]~q ),
	.datad(\Mux2~0_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hF388;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N2
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][29]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[18][29]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[26][29]~q ),
	.datad(\rfile[18][29]~q ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hB9A8;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y36_N8
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (instruction_D[23] & ((\Mux2~2_combout  & ((\rfile[30][29]~q ))) # (!\Mux2~2_combout  & (\rfile[22][29]~q )))) # (!instruction_D[23] & (((\Mux2~2_combout ))))

	.dataa(\rfile[22][29]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[30][29]~q ),
	.datad(\Mux2~2_combout ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'hF388;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y32_N1
dffeas \rfile[24][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][29] .is_wysiwyg = "true";
defparam \rfile[24][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X74_Y32_N23
dffeas \rfile[16][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][29] .is_wysiwyg = "true";
defparam \rfile[16][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N0
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[24][29]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[16][29]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[24][29]~q ),
	.datad(\rfile[16][29]~q ),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hB9A8;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N30
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (instruction_D[23] & ((\Mux2~4_combout  & (\rfile[28][29]~q )) # (!\Mux2~4_combout  & ((\rfile[20][29]~q ))))) # (!instruction_D[23] & (((\Mux2~4_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[28][29]~q ),
	.datac(\rfile[20][29]~q ),
	.datad(\Mux2~4_combout ),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hDDA0;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N28
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux2~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & ((\Mux2~5_combout ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux2~3_combout ),
	.datad(\Mux2~5_combout ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'hB9A8;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N14
cycloneive_lcell_comb \Mux2~17 (
// Equation(s):
// \Mux2~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][29]~q )) # (!instruction_D[21] & ((\rfile[12][29]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[13][29]~q ),
	.datad(\rfile[12][29]~q ),
	.cin(gnd),
	.combout(\Mux2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~17 .lut_mask = 16'hD9C8;
defparam \Mux2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N28
cycloneive_lcell_comb \Mux2~18 (
// Equation(s):
// \Mux2~18_combout  = (\Mux2~17_combout  & ((\rfile[15][29]~q ) # ((!instruction_D[22])))) # (!\Mux2~17_combout  & (((\rfile[14][29]~q  & instruction_D[22]))))

	.dataa(\Mux2~17_combout ),
	.datab(\rfile[15][29]~q ),
	.datac(\rfile[14][29]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~18 .lut_mask = 16'hD8AA;
defparam \Mux2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N10
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][29]~q )))) # (!instruction_D[22] & (!instruction_D[21] & (\rfile[8][29]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[8][29]~q ),
	.datad(\rfile[10][29]~q ),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'hBA98;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N4
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// \Mux2~11_combout  = (instruction_D[21] & ((\Mux2~10_combout  & ((\rfile[11][29]~q ))) # (!\Mux2~10_combout  & (\rfile[9][29]~q )))) # (!instruction_D[21] & (((\Mux2~10_combout ))))

	.dataa(\rfile[9][29]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[11][29]~q ),
	.datad(\Mux2~10_combout ),
	.cin(gnd),
	.combout(\Mux2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hF388;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N23
dffeas \rfile[7][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[7][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[7][29] .is_wysiwyg = "true";
defparam \rfile[7][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N24
cycloneive_lcell_comb \Mux2~12 (
// Equation(s):
// \Mux2~12_combout  = (instruction_D[21] & ((instruction_D[22]) # ((\rfile[5][29]~q )))) # (!instruction_D[21] & (!instruction_D[22] & ((\rfile[4][29]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[5][29]~q ),
	.datad(\rfile[4][29]~q ),
	.cin(gnd),
	.combout(\Mux2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~12 .lut_mask = 16'hB9A8;
defparam \Mux2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N22
cycloneive_lcell_comb \Mux2~13 (
// Equation(s):
// \Mux2~13_combout  = (instruction_D[22] & ((\Mux2~12_combout  & ((\rfile[7][29]~q ))) # (!\Mux2~12_combout  & (\rfile[6][29]~q )))) # (!instruction_D[22] & (((\Mux2~12_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[6][29]~q ),
	.datac(\rfile[7][29]~q ),
	.datad(\Mux2~12_combout ),
	.cin(gnd),
	.combout(\Mux2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~13 .lut_mask = 16'hF588;
defparam \Mux2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N0
cycloneive_lcell_comb \Mux2~14 (
// Equation(s):
// \Mux2~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][29]~q )) # (!instruction_D[22] & ((\rfile[1][29]~q )))))

	.dataa(instruction_D_22),
	.datab(\rfile[3][29]~q ),
	.datac(instruction_D_21),
	.datad(\rfile[1][29]~q ),
	.cin(gnd),
	.combout(\Mux2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~14 .lut_mask = 16'hD080;
defparam \Mux2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N18
cycloneive_lcell_comb \Mux2~15 (
// Equation(s):
// \Mux2~15_combout  = (\Mux2~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][29]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[2][29]~q ),
	.datad(\Mux2~14_combout ),
	.cin(gnd),
	.combout(\Mux2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~15 .lut_mask = 16'hFF20;
defparam \Mux2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N12
cycloneive_lcell_comb \Mux2~16 (
// Equation(s):
// \Mux2~16_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\Mux2~13_combout )))) # (!instruction_D[23] & (!instruction_D[24] & ((\Mux2~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux2~13_combout ),
	.datad(\Mux2~15_combout ),
	.cin(gnd),
	.combout(\Mux2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~16 .lut_mask = 16'hB9A8;
defparam \Mux2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y35_N15
dffeas \rfile[18][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][30] .is_wysiwyg = "true";
defparam \rfile[18][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N20
cycloneive_lcell_comb \rfile[22][30]~feeder (
// Equation(s):
// \rfile[22][30]~feeder_combout  = \wdat_WB[30]~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_30),
	.cin(gnd),
	.combout(\rfile[22][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[22][30]~feeder .lut_mask = 16'hFF00;
defparam \rfile[22][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y35_N21
dffeas \rfile[22][30] (
	.clk(!CLK),
	.d(\rfile[22][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][30] .is_wysiwyg = "true";
defparam \rfile[22][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N14
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// \Mux1~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[22][30]~q ))) # (!instruction_D[23] & (\rfile[18][30]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][30]~q ),
	.datad(\rfile[22][30]~q ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'hDC98;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N10
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (instruction_D[24] & ((\Mux1~2_combout  & ((\rfile[30][30]~q ))) # (!\Mux1~2_combout  & (\rfile[26][30]~q )))) # (!instruction_D[24] & (((\Mux1~2_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[26][30]~q ),
	.datac(\rfile[30][30]~q ),
	.datad(\Mux1~2_combout ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hF588;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N10
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[20][30]~q ))) # (!instruction_D[23] & (\rfile[16][30]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[16][30]~q ),
	.datad(\rfile[20][30]~q ),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'hDC98;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N14
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (instruction_D[24] & ((\Mux1~4_combout  & (\rfile[28][30]~q )) # (!\Mux1~4_combout  & ((\rfile[24][30]~q ))))) # (!instruction_D[24] & (((\Mux1~4_combout ))))

	.dataa(\rfile[28][30]~q ),
	.datab(instruction_D_24),
	.datac(\Mux1~4_combout ),
	.datad(\rfile[24][30]~q ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'hBCB0;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N12
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux1~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & ((\Mux1~5_combout ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux1~3_combout ),
	.datad(\Mux1~5_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hB9A8;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N14
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// \Mux1~7_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[27][30]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[19][30]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[19][30]~q ),
	.datad(\rfile[27][30]~q ),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hBA98;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N30
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// \Mux1~8_combout  = (instruction_D[23] & ((\Mux1~7_combout  & ((\rfile[31][30]~q ))) # (!\Mux1~7_combout  & (\rfile[23][30]~q )))) # (!instruction_D[23] & (((\Mux1~7_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[23][30]~q ),
	.datac(\rfile[31][30]~q ),
	.datad(\Mux1~7_combout ),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'hF588;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N18
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[25][30]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[17][30]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[17][30]~q ),
	.datad(\rfile[25][30]~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hBA98;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N16
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (\Mux1~0_combout  & (((\rfile[29][30]~q )) # (!instruction_D[23]))) # (!\Mux1~0_combout  & (instruction_D[23] & (\rfile[21][30]~q )))

	.dataa(\Mux1~0_combout ),
	.datab(instruction_D_23),
	.datac(\rfile[21][30]~q ),
	.datad(\rfile[29][30]~q ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hEA62;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N24
cycloneive_lcell_comb \Mux1~17 (
// Equation(s):
// \Mux1~17_combout  = (instruction_D[21] & ((\rfile[13][30]~q ) # ((instruction_D[22])))) # (!instruction_D[21] & (((\rfile[12][30]~q  & !instruction_D[22]))))

	.dataa(\rfile[13][30]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[12][30]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~17 .lut_mask = 16'hCCB8;
defparam \Mux1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N0
cycloneive_lcell_comb \Mux1~18 (
// Equation(s):
// \Mux1~18_combout  = (instruction_D[22] & ((\Mux1~17_combout  & (\rfile[15][30]~q )) # (!\Mux1~17_combout  & ((\rfile[14][30]~q ))))) # (!instruction_D[22] & (((\Mux1~17_combout ))))

	.dataa(\rfile[15][30]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[14][30]~q ),
	.datad(\Mux1~17_combout ),
	.cin(gnd),
	.combout(\Mux1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~18 .lut_mask = 16'hBBC0;
defparam \Mux1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N23
dffeas \rfile[4][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][30] .is_wysiwyg = "true";
defparam \rfile[4][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N22
cycloneive_lcell_comb \Mux1~10 (
// Equation(s):
// \Mux1~10_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[5][30]~q )) # (!instruction_D[21] & ((\rfile[4][30]~q )))))

	.dataa(instruction_D_22),
	.datab(\rfile[5][30]~q ),
	.datac(\rfile[4][30]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~10 .lut_mask = 16'hEE50;
defparam \Mux1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N2
cycloneive_lcell_comb \Mux1~11 (
// Equation(s):
// \Mux1~11_combout  = (instruction_D[22] & ((\Mux1~10_combout  & ((\rfile[7][30]~q ))) # (!\Mux1~10_combout  & (\rfile[6][30]~q )))) # (!instruction_D[22] & (((\Mux1~10_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[6][30]~q ),
	.datac(\rfile[7][30]~q ),
	.datad(\Mux1~10_combout ),
	.cin(gnd),
	.combout(\Mux1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~11 .lut_mask = 16'hF588;
defparam \Mux1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N6
cycloneive_lcell_comb \Mux1~14 (
// Equation(s):
// \Mux1~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][30]~q ))) # (!instruction_D[22] & (\rfile[1][30]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][30]~q ),
	.datad(\rfile[3][30]~q ),
	.cin(gnd),
	.combout(\Mux1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~14 .lut_mask = 16'hC840;
defparam \Mux1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N8
cycloneive_lcell_comb \Mux1~15 (
// Equation(s):
// \Mux1~15_combout  = (\Mux1~14_combout ) # ((!instruction_D[21] & (\rfile[2][30]~q  & instruction_D[22])))

	.dataa(instruction_D_21),
	.datab(\Mux1~14_combout ),
	.datac(\rfile[2][30]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~15 .lut_mask = 16'hDCCC;
defparam \Mux1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N31
dffeas \rfile[11][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][30] .is_wysiwyg = "true";
defparam \rfile[11][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N24
cycloneive_lcell_comb \Mux1~12 (
// Equation(s):
// \Mux1~12_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][30]~q )))) # (!instruction_D[22] & (!instruction_D[21] & ((\rfile[8][30]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[10][30]~q ),
	.datad(\rfile[8][30]~q ),
	.cin(gnd),
	.combout(\Mux1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~12 .lut_mask = 16'hB9A8;
defparam \Mux1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N30
cycloneive_lcell_comb \Mux1~13 (
// Equation(s):
// \Mux1~13_combout  = (instruction_D[21] & ((\Mux1~12_combout  & ((\rfile[11][30]~q ))) # (!\Mux1~12_combout  & (\rfile[9][30]~q )))) # (!instruction_D[21] & (((\Mux1~12_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[9][30]~q ),
	.datac(\rfile[11][30]~q ),
	.datad(\Mux1~12_combout ),
	.cin(gnd),
	.combout(\Mux1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~13 .lut_mask = 16'hF588;
defparam \Mux1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N2
cycloneive_lcell_comb \Mux1~16 (
// Equation(s):
// \Mux1~16_combout  = (instruction_D[24] & (((instruction_D[23]) # (\Mux1~13_combout )))) # (!instruction_D[24] & (\Mux1~15_combout  & (!instruction_D[23])))

	.dataa(instruction_D_24),
	.datab(\Mux1~15_combout ),
	.datac(instruction_D_23),
	.datad(\Mux1~13_combout ),
	.cin(gnd),
	.combout(\Mux1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~16 .lut_mask = 16'hAEA4;
defparam \Mux1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N28
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (instruction_D[24] & (((\rfile[25][28]~q ) # (instruction_D[23])))) # (!instruction_D[24] & (\rfile[17][28]~q  & ((!instruction_D[23]))))

	.dataa(\rfile[17][28]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[25][28]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hCCE2;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N24
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (\Mux3~0_combout  & (((\rfile[29][28]~q )) # (!instruction_D[23]))) # (!\Mux3~0_combout  & (instruction_D[23] & ((\rfile[21][28]~q ))))

	.dataa(\Mux3~0_combout ),
	.datab(instruction_D_23),
	.datac(\rfile[29][28]~q ),
	.datad(\rfile[21][28]~q ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hE6A2;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N2
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// \Mux3~7_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[27][28]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[19][28]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[19][28]~q ),
	.datad(\rfile[27][28]~q ),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hBA98;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N10
cycloneive_lcell_comb \Mux3~8 (
// Equation(s):
// \Mux3~8_combout  = (instruction_D[23] & ((\Mux3~7_combout  & (\rfile[31][28]~q )) # (!\Mux3~7_combout  & ((\rfile[23][28]~q ))))) # (!instruction_D[23] & (\Mux3~7_combout ))

	.dataa(instruction_D_23),
	.datab(\Mux3~7_combout ),
	.datac(\rfile[31][28]~q ),
	.datad(\rfile[23][28]~q ),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~8 .lut_mask = 16'hE6C4;
defparam \Mux3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N16
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[22][28]~q )) # (!instruction_D[23] & ((\rfile[18][28]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[22][28]~q ),
	.datad(\rfile[18][28]~q ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hD9C8;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N20
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (instruction_D[24] & ((\Mux3~2_combout  & (\rfile[30][28]~q )) # (!\Mux3~2_combout  & ((\rfile[26][28]~q ))))) # (!instruction_D[24] & (((\Mux3~2_combout ))))

	.dataa(\rfile[30][28]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[26][28]~q ),
	.datad(\Mux3~2_combout ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hBBC0;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N23
dffeas \rfile[28][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][28] .is_wysiwyg = "true";
defparam \rfile[28][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N28
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[20][28]~q )) # (!instruction_D[23] & ((\rfile[16][28]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[20][28]~q ),
	.datad(\rfile[16][28]~q ),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'hD9C8;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N22
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (instruction_D[24] & ((\Mux3~4_combout  & ((\rfile[28][28]~q ))) # (!\Mux3~4_combout  & (\rfile[24][28]~q )))) # (!instruction_D[24] & (((\Mux3~4_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[24][28]~q ),
	.datac(\rfile[28][28]~q ),
	.datad(\Mux3~4_combout ),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'hF588;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N2
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux3~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & ((\Mux3~5_combout ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux3~3_combout ),
	.datad(\Mux3~5_combout ),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'hB9A8;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N20
cycloneive_lcell_comb \Mux3~10 (
// Equation(s):
// \Mux3~10_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[5][28]~q ))) # (!instruction_D[21] & (\rfile[4][28]~q ))))

	.dataa(instruction_D_22),
	.datab(\rfile[4][28]~q ),
	.datac(\rfile[5][28]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~10 .lut_mask = 16'hFA44;
defparam \Mux3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N20
cycloneive_lcell_comb \Mux3~11 (
// Equation(s):
// \Mux3~11_combout  = (instruction_D[22] & ((\Mux3~10_combout  & (\rfile[7][28]~q )) # (!\Mux3~10_combout  & ((\rfile[6][28]~q ))))) # (!instruction_D[22] & (((\Mux3~10_combout ))))

	.dataa(\rfile[7][28]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[6][28]~q ),
	.datad(\Mux3~10_combout ),
	.cin(gnd),
	.combout(\Mux3~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~11 .lut_mask = 16'hBBC0;
defparam \Mux3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N10
cycloneive_lcell_comb \Mux3~17 (
// Equation(s):
// \Mux3~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][28]~q ))) # (!instruction_D[21] & (\rfile[12][28]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][28]~q ),
	.datad(\rfile[13][28]~q ),
	.cin(gnd),
	.combout(\Mux3~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~17 .lut_mask = 16'hDC98;
defparam \Mux3~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N26
cycloneive_lcell_comb \Mux3~18 (
// Equation(s):
// \Mux3~18_combout  = (instruction_D[22] & ((\Mux3~17_combout  & ((\rfile[15][28]~q ))) # (!\Mux3~17_combout  & (\rfile[14][28]~q )))) # (!instruction_D[22] & (((\Mux3~17_combout ))))

	.dataa(\rfile[14][28]~q ),
	.datab(instruction_D_22),
	.datac(\Mux3~17_combout ),
	.datad(\rfile[15][28]~q ),
	.cin(gnd),
	.combout(\Mux3~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~18 .lut_mask = 16'hF838;
defparam \Mux3~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N18
cycloneive_lcell_comb \Mux3~14 (
// Equation(s):
// \Mux3~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][28]~q ))) # (!instruction_D[22] & (\rfile[1][28]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][28]~q ),
	.datad(\rfile[3][28]~q ),
	.cin(gnd),
	.combout(\Mux3~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~14 .lut_mask = 16'hC840;
defparam \Mux3~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N22
cycloneive_lcell_comb \Mux3~15 (
// Equation(s):
// \Mux3~15_combout  = (\Mux3~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][28]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[2][28]~q ),
	.datad(\Mux3~14_combout ),
	.cin(gnd),
	.combout(\Mux3~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~15 .lut_mask = 16'hFF20;
defparam \Mux3~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N12
cycloneive_lcell_comb \Mux3~12 (
// Equation(s):
// \Mux3~12_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][28]~q )))) # (!instruction_D[22] & (!instruction_D[21] & ((\rfile[8][28]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[10][28]~q ),
	.datad(\rfile[8][28]~q ),
	.cin(gnd),
	.combout(\Mux3~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~12 .lut_mask = 16'hB9A8;
defparam \Mux3~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N6
cycloneive_lcell_comb \Mux3~13 (
// Equation(s):
// \Mux3~13_combout  = (instruction_D[21] & ((\Mux3~12_combout  & ((\rfile[11][28]~q ))) # (!\Mux3~12_combout  & (\rfile[9][28]~q )))) # (!instruction_D[21] & (((\Mux3~12_combout ))))

	.dataa(\rfile[9][28]~q ),
	.datab(\rfile[11][28]~q ),
	.datac(instruction_D_21),
	.datad(\Mux3~12_combout ),
	.cin(gnd),
	.combout(\Mux3~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~13 .lut_mask = 16'hCFA0;
defparam \Mux3~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N4
cycloneive_lcell_comb \Mux3~16 (
// Equation(s):
// \Mux3~16_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\Mux3~13_combout ))) # (!instruction_D[24] & (\Mux3~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux3~15_combout ),
	.datad(\Mux3~13_combout ),
	.cin(gnd),
	.combout(\Mux3~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~16 .lut_mask = 16'hDC98;
defparam \Mux3~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N8
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[21][27]~q )))) # (!instruction_D[23] & (!instruction_D[24] & ((\rfile[17][27]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[21][27]~q ),
	.datad(\rfile[17][27]~q ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hB9A8;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N14
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (\Mux4~0_combout  & (((\rfile[29][27]~q ) # (!instruction_D[24])))) # (!\Mux4~0_combout  & (\rfile[25][27]~q  & ((instruction_D[24]))))

	.dataa(\rfile[25][27]~q ),
	.datab(\rfile[29][27]~q ),
	.datac(\Mux4~0_combout ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hCAF0;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y29_N31
dffeas \rfile[19][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][27] .is_wysiwyg = "true";
defparam \rfile[19][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N30
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// \Mux4~7_combout  = (instruction_D[24] & (((instruction_D[23])))) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[23][27]~q )) # (!instruction_D[23] & ((\rfile[19][27]~q )))))

	.dataa(instruction_D_24),
	.datab(\rfile[23][27]~q ),
	.datac(\rfile[19][27]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'hEE50;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N18
cycloneive_lcell_comb \Mux4~8 (
// Equation(s):
// \Mux4~8_combout  = (\Mux4~7_combout  & (((\rfile[31][27]~q ) # (!instruction_D[24])))) # (!\Mux4~7_combout  & (\rfile[27][27]~q  & ((instruction_D[24]))))

	.dataa(\Mux4~7_combout ),
	.datab(\rfile[27][27]~q ),
	.datac(\rfile[31][27]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~8 .lut_mask = 16'hE4AA;
defparam \Mux4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N17
dffeas \rfile[22][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][27] .is_wysiwyg = "true";
defparam \rfile[22][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N18
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][27]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[18][27]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][27]~q ),
	.datad(\rfile[26][27]~q ),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hBA98;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N16
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (instruction_D[23] & ((\Mux4~2_combout  & (\rfile[30][27]~q )) # (!\Mux4~2_combout  & ((\rfile[22][27]~q ))))) # (!instruction_D[23] & (((\Mux4~2_combout ))))

	.dataa(\rfile[30][27]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[22][27]~q ),
	.datad(\Mux4~2_combout ),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hBBC0;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N5
dffeas \rfile[28][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][27] .is_wysiwyg = "true";
defparam \rfile[28][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y32_N16
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[24][27]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[16][27]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[16][27]~q ),
	.datad(\rfile[24][27]~q ),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'hBA98;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N4
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (instruction_D[23] & ((\Mux4~4_combout  & ((\rfile[28][27]~q ))) # (!\Mux4~4_combout  & (\rfile[20][27]~q )))) # (!instruction_D[23] & (((\Mux4~4_combout ))))

	.dataa(\rfile[20][27]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[28][27]~q ),
	.datad(\Mux4~4_combout ),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'hF388;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N16
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// \Mux4~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux4~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & ((\Mux4~5_combout ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux4~3_combout ),
	.datad(\Mux4~5_combout ),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hB9A8;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N6
cycloneive_lcell_comb \Mux4~17 (
// Equation(s):
// \Mux4~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][27]~q ))) # (!instruction_D[21] & (\rfile[12][27]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][27]~q ),
	.datad(\rfile[13][27]~q ),
	.cin(gnd),
	.combout(\Mux4~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~17 .lut_mask = 16'hDC98;
defparam \Mux4~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N16
cycloneive_lcell_comb \Mux4~18 (
// Equation(s):
// \Mux4~18_combout  = (\Mux4~17_combout  & (((\rfile[15][27]~q ) # (!instruction_D[22])))) # (!\Mux4~17_combout  & (\rfile[14][27]~q  & ((instruction_D[22]))))

	.dataa(\rfile[14][27]~q ),
	.datab(\Mux4~17_combout ),
	.datac(\rfile[15][27]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux4~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~18 .lut_mask = 16'hE2CC;
defparam \Mux4~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N16
cycloneive_lcell_comb \Mux4~10 (
// Equation(s):
// \Mux4~10_combout  = (instruction_D[21] & (((instruction_D[22])))) # (!instruction_D[21] & ((instruction_D[22] & ((\rfile[10][27]~q ))) # (!instruction_D[22] & (\rfile[8][27]~q ))))

	.dataa(\rfile[8][27]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[10][27]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux4~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~10 .lut_mask = 16'hFC22;
defparam \Mux4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N20
cycloneive_lcell_comb \Mux4~11 (
// Equation(s):
// \Mux4~11_combout  = (instruction_D[21] & ((\Mux4~10_combout  & (\rfile[11][27]~q )) # (!\Mux4~10_combout  & ((\rfile[9][27]~q ))))) # (!instruction_D[21] & (((\Mux4~10_combout ))))

	.dataa(\rfile[11][27]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[9][27]~q ),
	.datad(\Mux4~10_combout ),
	.cin(gnd),
	.combout(\Mux4~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~11 .lut_mask = 16'hBBC0;
defparam \Mux4~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N22
cycloneive_lcell_comb \Mux4~14 (
// Equation(s):
// \Mux4~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][27]~q ))) # (!instruction_D[22] & (\rfile[1][27]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][27]~q ),
	.datad(\rfile[3][27]~q ),
	.cin(gnd),
	.combout(\Mux4~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~14 .lut_mask = 16'hC840;
defparam \Mux4~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N30
cycloneive_lcell_comb \Mux4~15 (
// Equation(s):
// \Mux4~15_combout  = (\Mux4~14_combout ) # ((instruction_D[22] & (\rfile[2][27]~q  & !instruction_D[21])))

	.dataa(instruction_D_22),
	.datab(\rfile[2][27]~q ),
	.datac(instruction_D_21),
	.datad(\Mux4~14_combout ),
	.cin(gnd),
	.combout(\Mux4~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~15 .lut_mask = 16'hFF08;
defparam \Mux4~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N10
cycloneive_lcell_comb \Mux4~12 (
// Equation(s):
// \Mux4~12_combout  = (instruction_D[21] & ((instruction_D[22]) # ((\rfile[5][27]~q )))) # (!instruction_D[21] & (!instruction_D[22] & (\rfile[4][27]~q )))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[4][27]~q ),
	.datad(\rfile[5][27]~q ),
	.cin(gnd),
	.combout(\Mux4~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~12 .lut_mask = 16'hBA98;
defparam \Mux4~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N10
cycloneive_lcell_comb \Mux4~13 (
// Equation(s):
// \Mux4~13_combout  = (instruction_D[22] & ((\Mux4~12_combout  & (\rfile[7][27]~q )) # (!\Mux4~12_combout  & ((\rfile[6][27]~q ))))) # (!instruction_D[22] & (((\Mux4~12_combout ))))

	.dataa(\rfile[7][27]~q ),
	.datab(\rfile[6][27]~q ),
	.datac(instruction_D_22),
	.datad(\Mux4~12_combout ),
	.cin(gnd),
	.combout(\Mux4~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~13 .lut_mask = 16'hAFC0;
defparam \Mux4~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N12
cycloneive_lcell_comb \Mux4~16 (
// Equation(s):
// \Mux4~16_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\Mux4~13_combout )))) # (!instruction_D[23] & (!instruction_D[24] & (\Mux4~15_combout )))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux4~15_combout ),
	.datad(\Mux4~13_combout ),
	.cin(gnd),
	.combout(\Mux4~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~16 .lut_mask = 16'hBA98;
defparam \Mux4~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y27_N27
dffeas \rfile[17][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[17][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[17][26] .is_wysiwyg = "true";
defparam \rfile[17][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N26
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[25][26]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[17][26]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[17][26]~q ),
	.datad(\rfile[25][26]~q ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hBA98;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N30
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (instruction_D[23] & ((\Mux5~0_combout  & ((\rfile[29][26]~q ))) # (!\Mux5~0_combout  & (\rfile[21][26]~q )))) # (!instruction_D[23] & (\Mux5~0_combout ))

	.dataa(instruction_D_23),
	.datab(\Mux5~0_combout ),
	.datac(\rfile[21][26]~q ),
	.datad(\rfile[29][26]~q ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hEC64;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N10
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[27][26]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[19][26]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[19][26]~q ),
	.datad(\rfile[27][26]~q ),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'hBA98;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N26
cycloneive_lcell_comb \Mux5~8 (
// Equation(s):
// \Mux5~8_combout  = (instruction_D[23] & ((\Mux5~7_combout  & (\rfile[31][26]~q )) # (!\Mux5~7_combout  & ((\rfile[23][26]~q ))))) # (!instruction_D[23] & (((\Mux5~7_combout ))))

	.dataa(\rfile[31][26]~q ),
	.datab(instruction_D_23),
	.datac(\Mux5~7_combout ),
	.datad(\rfile[23][26]~q ),
	.cin(gnd),
	.combout(\Mux5~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~8 .lut_mask = 16'hBCB0;
defparam \Mux5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y31_N27
dffeas \rfile[16][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[16][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[16][26] .is_wysiwyg = "true";
defparam \rfile[16][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X76_Y31_N21
dffeas \rfile[20][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][26] .is_wysiwyg = "true";
defparam \rfile[20][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N26
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[20][26]~q ))) # (!instruction_D[23] & (\rfile[16][26]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[16][26]~q ),
	.datad(\rfile[20][26]~q ),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'hDC98;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N6
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (instruction_D[24] & ((\Mux5~4_combout  & ((\rfile[28][26]~q ))) # (!\Mux5~4_combout  & (\rfile[24][26]~q )))) # (!instruction_D[24] & (((\Mux5~4_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[24][26]~q ),
	.datac(\rfile[28][26]~q ),
	.datad(\Mux5~4_combout ),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'hF588;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y34_N31
dffeas \rfile[18][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][26] .is_wysiwyg = "true";
defparam \rfile[18][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N30
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (instruction_D[24] & (((instruction_D[23])))) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[22][26]~q )) # (!instruction_D[23] & ((\rfile[18][26]~q )))))

	.dataa(instruction_D_24),
	.datab(\rfile[22][26]~q ),
	.datac(\rfile[18][26]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hEE50;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N2
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (instruction_D[24] & ((\Mux5~2_combout  & ((\rfile[30][26]~q ))) # (!\Mux5~2_combout  & (\rfile[26][26]~q )))) # (!instruction_D[24] & (((\Mux5~2_combout ))))

	.dataa(\rfile[26][26]~q ),
	.datab(instruction_D_24),
	.datac(\Mux5~2_combout ),
	.datad(\rfile[30][26]~q ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hF838;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N26
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux5~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & (\Mux5~5_combout )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux5~5_combout ),
	.datad(\Mux5~3_combout ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hBA98;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N16
cycloneive_lcell_comb \Mux5~10 (
// Equation(s):
// \Mux5~10_combout  = (instruction_D[21] & ((instruction_D[22]) # ((\rfile[5][26]~q )))) # (!instruction_D[21] & (!instruction_D[22] & ((\rfile[4][26]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[5][26]~q ),
	.datad(\rfile[4][26]~q ),
	.cin(gnd),
	.combout(\Mux5~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~10 .lut_mask = 16'hB9A8;
defparam \Mux5~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N12
cycloneive_lcell_comb \Mux5~11 (
// Equation(s):
// \Mux5~11_combout  = (instruction_D[22] & ((\Mux5~10_combout  & (\rfile[7][26]~q )) # (!\Mux5~10_combout  & ((\rfile[6][26]~q ))))) # (!instruction_D[22] & (((\Mux5~10_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[7][26]~q ),
	.datac(\rfile[6][26]~q ),
	.datad(\Mux5~10_combout ),
	.cin(gnd),
	.combout(\Mux5~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~11 .lut_mask = 16'hDDA0;
defparam \Mux5~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N20
cycloneive_lcell_comb \Mux5~17 (
// Equation(s):
// \Mux5~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][26]~q )) # (!instruction_D[21] & ((\rfile[12][26]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[13][26]~q ),
	.datad(\rfile[12][26]~q ),
	.cin(gnd),
	.combout(\Mux5~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~17 .lut_mask = 16'hD9C8;
defparam \Mux5~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N24
cycloneive_lcell_comb \Mux5~18 (
// Equation(s):
// \Mux5~18_combout  = (instruction_D[22] & ((\Mux5~17_combout  & ((\rfile[15][26]~q ))) # (!\Mux5~17_combout  & (\rfile[14][26]~q )))) # (!instruction_D[22] & (((\Mux5~17_combout ))))

	.dataa(\rfile[14][26]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[15][26]~q ),
	.datad(\Mux5~17_combout ),
	.cin(gnd),
	.combout(\Mux5~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~18 .lut_mask = 16'hF388;
defparam \Mux5~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N24
cycloneive_lcell_comb \Mux5~14 (
// Equation(s):
// \Mux5~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][26]~q )) # (!instruction_D[22] & ((\rfile[1][26]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[3][26]~q ),
	.datad(\rfile[1][26]~q ),
	.cin(gnd),
	.combout(\Mux5~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~14 .lut_mask = 16'hC480;
defparam \Mux5~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N26
cycloneive_lcell_comb \Mux5~15 (
// Equation(s):
// \Mux5~15_combout  = (\Mux5~14_combout ) # ((\rfile[2][26]~q  & (!instruction_D[21] & instruction_D[22])))

	.dataa(\rfile[2][26]~q ),
	.datab(instruction_D_21),
	.datac(instruction_D_22),
	.datad(\Mux5~14_combout ),
	.cin(gnd),
	.combout(\Mux5~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~15 .lut_mask = 16'hFF20;
defparam \Mux5~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N17
dffeas \rfile[11][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][26] .is_wysiwyg = "true";
defparam \rfile[11][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N9
dffeas \rfile[10][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[10][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[10][26] .is_wysiwyg = "true";
defparam \rfile[10][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N8
cycloneive_lcell_comb \Mux5~12 (
// Equation(s):
// \Mux5~12_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][26]~q )))) # (!instruction_D[22] & (!instruction_D[21] & ((\rfile[8][26]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[10][26]~q ),
	.datad(\rfile[8][26]~q ),
	.cin(gnd),
	.combout(\Mux5~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~12 .lut_mask = 16'hB9A8;
defparam \Mux5~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N16
cycloneive_lcell_comb \Mux5~13 (
// Equation(s):
// \Mux5~13_combout  = (instruction_D[21] & ((\Mux5~12_combout  & ((\rfile[11][26]~q ))) # (!\Mux5~12_combout  & (\rfile[9][26]~q )))) # (!instruction_D[21] & (((\Mux5~12_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[9][26]~q ),
	.datac(\rfile[11][26]~q ),
	.datad(\Mux5~12_combout ),
	.cin(gnd),
	.combout(\Mux5~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~13 .lut_mask = 16'hF588;
defparam \Mux5~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N28
cycloneive_lcell_comb \Mux5~16 (
// Equation(s):
// \Mux5~16_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\Mux5~13_combout )))) # (!instruction_D[24] & (!instruction_D[23] & (\Mux5~15_combout )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux5~15_combout ),
	.datad(\Mux5~13_combout ),
	.cin(gnd),
	.combout(\Mux5~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~16 .lut_mask = 16'hBA98;
defparam \Mux5~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y29_N23
dffeas \rfile[19][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[19][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[19][25] .is_wysiwyg = "true";
defparam \rfile[19][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N22
cycloneive_lcell_comb \Mux6~7 (
// Equation(s):
// \Mux6~7_combout  = (instruction_D[24] & (((instruction_D[23])))) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[23][25]~q )) # (!instruction_D[23] & ((\rfile[19][25]~q )))))

	.dataa(instruction_D_24),
	.datab(\rfile[23][25]~q ),
	.datac(\rfile[19][25]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~7 .lut_mask = 16'hEE50;
defparam \Mux6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N14
cycloneive_lcell_comb \Mux6~8 (
// Equation(s):
// \Mux6~8_combout  = (instruction_D[24] & ((\Mux6~7_combout  & ((\rfile[31][25]~q ))) # (!\Mux6~7_combout  & (\rfile[27][25]~q )))) # (!instruction_D[24] & (((\Mux6~7_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[27][25]~q ),
	.datac(\rfile[31][25]~q ),
	.datad(\Mux6~7_combout ),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~8 .lut_mask = 16'hF588;
defparam \Mux6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N0
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[21][25]~q ))) # (!instruction_D[23] & (\rfile[17][25]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[17][25]~q ),
	.datad(\rfile[21][25]~q ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hDC98;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N14
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (instruction_D[24] & ((\Mux6~0_combout  & ((\rfile[29][25]~q ))) # (!\Mux6~0_combout  & (\rfile[25][25]~q )))) # (!instruction_D[24] & (((\Mux6~0_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[25][25]~q ),
	.datac(\rfile[29][25]~q ),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hF588;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y35_N23
dffeas \rfile[18][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[18][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[18][25] .is_wysiwyg = "true";
defparam \rfile[18][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N1
dffeas \rfile[26][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[26][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[26][25] .is_wysiwyg = "true";
defparam \rfile[26][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N22
cycloneive_lcell_comb \Mux6~2 (
// Equation(s):
// \Mux6~2_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\rfile[26][25]~q ))) # (!instruction_D[24] & (\rfile[18][25]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[18][25]~q ),
	.datad(\rfile[26][25]~q ),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~2 .lut_mask = 16'hDC98;
defparam \Mux6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N28
cycloneive_lcell_comb \Mux6~3 (
// Equation(s):
// \Mux6~3_combout  = (instruction_D[23] & ((\Mux6~2_combout  & (\rfile[30][25]~q )) # (!\Mux6~2_combout  & ((\rfile[22][25]~q ))))) # (!instruction_D[23] & (((\Mux6~2_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[30][25]~q ),
	.datac(\rfile[22][25]~q ),
	.datad(\Mux6~2_combout ),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~3 .lut_mask = 16'hDDA0;
defparam \Mux6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y31_N4
cycloneive_lcell_comb \rfile[28][25]~feeder (
// Equation(s):
// \rfile[28][25]~feeder_combout  = \wdat_WB[25]~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_25),
	.cin(gnd),
	.combout(\rfile[28][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[28][25]~feeder .lut_mask = 16'hFF00;
defparam \rfile[28][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X77_Y31_N5
dffeas \rfile[28][25] (
	.clk(!CLK),
	.d(\rfile[28][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][25] .is_wysiwyg = "true";
defparam \rfile[28][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X77_Y32_N30
cycloneive_lcell_comb \Mux6~4 (
// Equation(s):
// \Mux6~4_combout  = (instruction_D[23] & (((instruction_D[24])))) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[24][25]~q )) # (!instruction_D[24] & ((\rfile[16][25]~q )))))

	.dataa(\rfile[24][25]~q ),
	.datab(instruction_D_23),
	.datac(instruction_D_24),
	.datad(\rfile[16][25]~q ),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~4 .lut_mask = 16'hE3E0;
defparam \Mux6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X77_Y31_N2
cycloneive_lcell_comb \Mux6~5 (
// Equation(s):
// \Mux6~5_combout  = (instruction_D[23] & ((\Mux6~4_combout  & (\rfile[28][25]~q )) # (!\Mux6~4_combout  & ((\rfile[20][25]~q ))))) # (!instruction_D[23] & (((\Mux6~4_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[28][25]~q ),
	.datac(\Mux6~4_combout ),
	.datad(\rfile[20][25]~q ),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~5 .lut_mask = 16'hDAD0;
defparam \Mux6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N18
cycloneive_lcell_comb \Mux6~6 (
// Equation(s):
// \Mux6~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux6~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & ((\Mux6~5_combout ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux6~3_combout ),
	.datad(\Mux6~5_combout ),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~6 .lut_mask = 16'hB9A8;
defparam \Mux6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N4
cycloneive_lcell_comb \Mux6~10 (
// Equation(s):
// \Mux6~10_combout  = (instruction_D[21] & (((instruction_D[22])))) # (!instruction_D[21] & ((instruction_D[22] & ((\rfile[10][25]~q ))) # (!instruction_D[22] & (\rfile[8][25]~q ))))

	.dataa(\rfile[8][25]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[10][25]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux6~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~10 .lut_mask = 16'hFC22;
defparam \Mux6~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N12
cycloneive_lcell_comb \Mux6~11 (
// Equation(s):
// \Mux6~11_combout  = (instruction_D[21] & ((\Mux6~10_combout  & (\rfile[11][25]~q )) # (!\Mux6~10_combout  & ((\rfile[9][25]~q ))))) # (!instruction_D[21] & (((\Mux6~10_combout ))))

	.dataa(\rfile[11][25]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[9][25]~q ),
	.datad(\Mux6~10_combout ),
	.cin(gnd),
	.combout(\Mux6~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~11 .lut_mask = 16'hBBC0;
defparam \Mux6~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N18
cycloneive_lcell_comb \Mux6~14 (
// Equation(s):
// \Mux6~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][25]~q )) # (!instruction_D[22] & ((\rfile[1][25]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[3][25]~q ),
	.datad(\rfile[1][25]~q ),
	.cin(gnd),
	.combout(\Mux6~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~14 .lut_mask = 16'hC480;
defparam \Mux6~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N22
cycloneive_lcell_comb \Mux6~15 (
// Equation(s):
// \Mux6~15_combout  = (\Mux6~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][25]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[2][25]~q ),
	.datad(\Mux6~14_combout ),
	.cin(gnd),
	.combout(\Mux6~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~15 .lut_mask = 16'hFF20;
defparam \Mux6~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N2
cycloneive_lcell_comb \Mux6~12 (
// Equation(s):
// \Mux6~12_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[5][25]~q )) # (!instruction_D[21] & ((\rfile[4][25]~q )))))

	.dataa(instruction_D_22),
	.datab(\rfile[5][25]~q ),
	.datac(\rfile[4][25]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux6~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~12 .lut_mask = 16'hEE50;
defparam \Mux6~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N14
cycloneive_lcell_comb \Mux6~13 (
// Equation(s):
// \Mux6~13_combout  = (instruction_D[22] & ((\Mux6~12_combout  & ((\rfile[7][25]~q ))) # (!\Mux6~12_combout  & (\rfile[6][25]~q )))) # (!instruction_D[22] & (((\Mux6~12_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[6][25]~q ),
	.datac(\rfile[7][25]~q ),
	.datad(\Mux6~12_combout ),
	.cin(gnd),
	.combout(\Mux6~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~13 .lut_mask = 16'hF588;
defparam \Mux6~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N22
cycloneive_lcell_comb \Mux6~16 (
// Equation(s):
// \Mux6~16_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\Mux6~13_combout ))) # (!instruction_D[23] & (\Mux6~15_combout ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux6~15_combout ),
	.datad(\Mux6~13_combout ),
	.cin(gnd),
	.combout(\Mux6~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~16 .lut_mask = 16'hDC98;
defparam \Mux6~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N16
cycloneive_lcell_comb \Mux6~17 (
// Equation(s):
// \Mux6~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][25]~q )) # (!instruction_D[21] & ((\rfile[12][25]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[13][25]~q ),
	.datad(\rfile[12][25]~q ),
	.cin(gnd),
	.combout(\Mux6~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~17 .lut_mask = 16'hD9C8;
defparam \Mux6~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N4
cycloneive_lcell_comb \Mux6~18 (
// Equation(s):
// \Mux6~18_combout  = (instruction_D[22] & ((\Mux6~17_combout  & (\rfile[15][25]~q )) # (!\Mux6~17_combout  & ((\rfile[14][25]~q ))))) # (!instruction_D[22] & (((\Mux6~17_combout ))))

	.dataa(\rfile[15][25]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[14][25]~q ),
	.datad(\Mux6~17_combout ),
	.cin(gnd),
	.combout(\Mux6~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~18 .lut_mask = 16'hBBC0;
defparam \Mux6~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N4
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// \Mux7~7_combout  = (instruction_D[23] & (((instruction_D[24])))) # (!instruction_D[23] & ((instruction_D[24] & ((\rfile[27][24]~q ))) # (!instruction_D[24] & (\rfile[19][24]~q ))))

	.dataa(\rfile[19][24]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[27][24]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'hFC22;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N18
cycloneive_lcell_comb \Mux7~8 (
// Equation(s):
// \Mux7~8_combout  = (instruction_D[23] & ((\Mux7~7_combout  & (\rfile[31][24]~q )) # (!\Mux7~7_combout  & ((\rfile[23][24]~q ))))) # (!instruction_D[23] & (((\Mux7~7_combout ))))

	.dataa(\rfile[31][24]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[23][24]~q ),
	.datad(\Mux7~7_combout ),
	.cin(gnd),
	.combout(\Mux7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~8 .lut_mask = 16'hBBC0;
defparam \Mux7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N14
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[25][24]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[17][24]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[25][24]~q ),
	.datad(\rfile[17][24]~q ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hB9A8;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N14
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (instruction_D[23] & ((\Mux7~0_combout  & ((\rfile[29][24]~q ))) # (!\Mux7~0_combout  & (\rfile[21][24]~q )))) # (!instruction_D[23] & (((\Mux7~0_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[21][24]~q ),
	.datac(\rfile[29][24]~q ),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hF588;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N18
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (\Mux7~2_combout  & (((\rfile[30][24]~q )) # (!instruction_D[24]))) # (!\Mux7~2_combout  & (instruction_D[24] & (\rfile[26][24]~q )))

	.dataa(\Mux7~2_combout ),
	.datab(instruction_D_24),
	.datac(\rfile[26][24]~q ),
	.datad(\rfile[30][24]~q ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'hEA62;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X76_Y31_N5
dffeas \rfile[20][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][24] .is_wysiwyg = "true";
defparam \rfile[20][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N4
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (instruction_D[23] & (((\rfile[20][24]~q ) # (instruction_D[24])))) # (!instruction_D[23] & (\rfile[16][24]~q  & ((!instruction_D[24]))))

	.dataa(\rfile[16][24]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[20][24]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'hCCE2;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N28
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (instruction_D[24] & ((\Mux7~4_combout  & (\rfile[28][24]~q )) # (!\Mux7~4_combout  & ((\rfile[24][24]~q ))))) # (!instruction_D[24] & (((\Mux7~4_combout ))))

	.dataa(\rfile[28][24]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[24][24]~q ),
	.datad(\Mux7~4_combout ),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'hBBC0;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N12
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// \Mux7~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\Mux7~3_combout )) # (!instruction_D[22] & ((\Mux7~5_combout )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux7~3_combout ),
	.datad(\Mux7~5_combout ),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'hD9C8;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N13
dffeas \rfile[4][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][24] .is_wysiwyg = "true";
defparam \rfile[4][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N12
cycloneive_lcell_comb \Mux7~10 (
// Equation(s):
// \Mux7~10_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[5][24]~q )) # (!instruction_D[21] & ((\rfile[4][24]~q )))))

	.dataa(instruction_D_22),
	.datab(\rfile[5][24]~q ),
	.datac(\rfile[4][24]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~10 .lut_mask = 16'hEE50;
defparam \Mux7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N22
cycloneive_lcell_comb \Mux7~11 (
// Equation(s):
// \Mux7~11_combout  = (instruction_D[22] & ((\Mux7~10_combout  & ((\rfile[7][24]~q ))) # (!\Mux7~10_combout  & (\rfile[6][24]~q )))) # (!instruction_D[22] & (((\Mux7~10_combout ))))

	.dataa(\rfile[6][24]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[7][24]~q ),
	.datad(\Mux7~10_combout ),
	.cin(gnd),
	.combout(\Mux7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~11 .lut_mask = 16'hF388;
defparam \Mux7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N20
cycloneive_lcell_comb \Mux7~14 (
// Equation(s):
// \Mux7~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][24]~q )) # (!instruction_D[22] & ((\rfile[1][24]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[3][24]~q ),
	.datad(\rfile[1][24]~q ),
	.cin(gnd),
	.combout(\Mux7~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~14 .lut_mask = 16'hC480;
defparam \Mux7~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N22
cycloneive_lcell_comb \Mux7~15 (
// Equation(s):
// \Mux7~15_combout  = (\Mux7~14_combout ) # ((!instruction_D[21] & (\rfile[2][24]~q  & instruction_D[22])))

	.dataa(instruction_D_21),
	.datab(\rfile[2][24]~q ),
	.datac(instruction_D_22),
	.datad(\Mux7~14_combout ),
	.cin(gnd),
	.combout(\Mux7~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~15 .lut_mask = 16'hFF40;
defparam \Mux7~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N0
cycloneive_lcell_comb \Mux7~12 (
// Equation(s):
// \Mux7~12_combout  = (instruction_D[22] & (((\rfile[10][24]~q ) # (instruction_D[21])))) # (!instruction_D[22] & (\rfile[8][24]~q  & ((!instruction_D[21]))))

	.dataa(\rfile[8][24]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[10][24]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux7~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~12 .lut_mask = 16'hCCE2;
defparam \Mux7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N24
cycloneive_lcell_comb \Mux7~13 (
// Equation(s):
// \Mux7~13_combout  = (\Mux7~12_combout  & (((\rfile[11][24]~q ) # (!instruction_D[21])))) # (!\Mux7~12_combout  & (\rfile[9][24]~q  & ((instruction_D[21]))))

	.dataa(\rfile[9][24]~q ),
	.datab(\rfile[11][24]~q ),
	.datac(\Mux7~12_combout ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~13 .lut_mask = 16'hCAF0;
defparam \Mux7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N4
cycloneive_lcell_comb \Mux7~16 (
// Equation(s):
// \Mux7~16_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\Mux7~13_combout )))) # (!instruction_D[24] & (!instruction_D[23] & (\Mux7~15_combout )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux7~15_combout ),
	.datad(\Mux7~13_combout ),
	.cin(gnd),
	.combout(\Mux7~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~16 .lut_mask = 16'hBA98;
defparam \Mux7~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N26
cycloneive_lcell_comb \Mux7~17 (
// Equation(s):
// \Mux7~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][24]~q ))) # (!instruction_D[21] & (\rfile[12][24]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][24]~q ),
	.datad(\rfile[13][24]~q ),
	.cin(gnd),
	.combout(\Mux7~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~17 .lut_mask = 16'hDC98;
defparam \Mux7~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N2
cycloneive_lcell_comb \Mux7~18 (
// Equation(s):
// \Mux7~18_combout  = (instruction_D[22] & ((\Mux7~17_combout  & ((\rfile[15][24]~q ))) # (!\Mux7~17_combout  & (\rfile[14][24]~q )))) # (!instruction_D[22] & (((\Mux7~17_combout ))))

	.dataa(\rfile[14][24]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[15][24]~q ),
	.datad(\Mux7~17_combout ),
	.cin(gnd),
	.combout(\Mux7~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~18 .lut_mask = 16'hF388;
defparam \Mux7~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N4
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[21][23]~q )))) # (!instruction_D[23] & (!instruction_D[24] & ((\rfile[17][23]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[21][23]~q ),
	.datad(\rfile[17][23]~q ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hB9A8;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N24
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (\Mux8~0_combout  & ((\rfile[29][23]~q ) # ((!instruction_D[24])))) # (!\Mux8~0_combout  & (((\rfile[25][23]~q  & instruction_D[24]))))

	.dataa(\Mux8~0_combout ),
	.datab(\rfile[29][23]~q ),
	.datac(\rfile[25][23]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hD8AA;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N12
cycloneive_lcell_comb \Mux8~7 (
// Equation(s):
// \Mux8~7_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[23][23]~q )) # (!instruction_D[23] & ((\rfile[19][23]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[23][23]~q ),
	.datad(\rfile[19][23]~q ),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~7 .lut_mask = 16'hD9C8;
defparam \Mux8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N28
cycloneive_lcell_comb \Mux8~8 (
// Equation(s):
// \Mux8~8_combout  = (instruction_D[24] & ((\Mux8~7_combout  & (\rfile[31][23]~q )) # (!\Mux8~7_combout  & ((\rfile[27][23]~q ))))) # (!instruction_D[24] & (((\Mux8~7_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[31][23]~q ),
	.datac(\rfile[27][23]~q ),
	.datad(\Mux8~7_combout ),
	.cin(gnd),
	.combout(\Mux8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~8 .lut_mask = 16'hDDA0;
defparam \Mux8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y32_N12
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[24][23]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[16][23]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[24][23]~q ),
	.datad(\rfile[16][23]~q ),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'hB9A8;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N24
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// \Mux8~5_combout  = (instruction_D[23] & ((\Mux8~4_combout  & (\rfile[28][23]~q )) # (!\Mux8~4_combout  & ((\rfile[20][23]~q ))))) # (!instruction_D[23] & (((\Mux8~4_combout ))))

	.dataa(\rfile[28][23]~q ),
	.datab(instruction_D_23),
	.datac(\Mux8~4_combout ),
	.datad(\rfile[20][23]~q ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'hBCB0;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y36_N12
cycloneive_lcell_comb \Mux8~2 (
// Equation(s):
// \Mux8~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][23]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[18][23]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][23]~q ),
	.datad(\rfile[26][23]~q ),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~2 .lut_mask = 16'hBA98;
defparam \Mux8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N26
cycloneive_lcell_comb \Mux8~3 (
// Equation(s):
// \Mux8~3_combout  = (instruction_D[23] & ((\Mux8~2_combout  & ((\rfile[30][23]~q ))) # (!\Mux8~2_combout  & (\rfile[22][23]~q )))) # (!instruction_D[23] & (((\Mux8~2_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[22][23]~q ),
	.datac(\rfile[30][23]~q ),
	.datad(\Mux8~2_combout ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~3 .lut_mask = 16'hF588;
defparam \Mux8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N28
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux8~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & (\Mux8~5_combout )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux8~5_combout ),
	.datad(\Mux8~3_combout ),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hBA98;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N2
cycloneive_lcell_comb \Mux8~17 (
// Equation(s):
// \Mux8~17_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[13][23]~q )) # (!instruction_D[21] & ((\rfile[12][23]~q )))))

	.dataa(instruction_D_22),
	.datab(\rfile[13][23]~q ),
	.datac(\rfile[12][23]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux8~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~17 .lut_mask = 16'hEE50;
defparam \Mux8~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N16
cycloneive_lcell_comb \Mux8~18 (
// Equation(s):
// \Mux8~18_combout  = (instruction_D[22] & ((\Mux8~17_combout  & (\rfile[15][23]~q )) # (!\Mux8~17_combout  & ((\rfile[14][23]~q ))))) # (!instruction_D[22] & (((\Mux8~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[15][23]~q ),
	.datac(\rfile[14][23]~q ),
	.datad(\Mux8~17_combout ),
	.cin(gnd),
	.combout(\Mux8~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~18 .lut_mask = 16'hDDA0;
defparam \Mux8~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N18
cycloneive_lcell_comb \Mux8~14 (
// Equation(s):
// \Mux8~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][23]~q ))) # (!instruction_D[22] & (\rfile[1][23]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][23]~q ),
	.datad(\rfile[3][23]~q ),
	.cin(gnd),
	.combout(\Mux8~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~14 .lut_mask = 16'hC840;
defparam \Mux8~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N4
cycloneive_lcell_comb \Mux8~15 (
// Equation(s):
// \Mux8~15_combout  = (\Mux8~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][23]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux8~14_combout ),
	.datad(\rfile[2][23]~q ),
	.cin(gnd),
	.combout(\Mux8~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~15 .lut_mask = 16'hF2F0;
defparam \Mux8~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N24
cycloneive_lcell_comb \Mux8~12 (
// Equation(s):
// \Mux8~12_combout  = (instruction_D[21] & ((\rfile[5][23]~q ) # ((instruction_D[22])))) # (!instruction_D[21] & (((\rfile[4][23]~q  & !instruction_D[22]))))

	.dataa(instruction_D_21),
	.datab(\rfile[5][23]~q ),
	.datac(\rfile[4][23]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux8~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~12 .lut_mask = 16'hAAD8;
defparam \Mux8~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N16
cycloneive_lcell_comb \rfile[6][23]~feeder (
// Equation(s):
// \rfile[6][23]~feeder_combout  = \wdat_WB[23]~19_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat_WB_23),
	.cin(gnd),
	.combout(\rfile[6][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[6][23]~feeder .lut_mask = 16'hFF00;
defparam \rfile[6][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N17
dffeas \rfile[6][23] (
	.clk(!CLK),
	.d(\rfile[6][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[6][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[6][23] .is_wysiwyg = "true";
defparam \rfile[6][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N2
cycloneive_lcell_comb \Mux8~13 (
// Equation(s):
// \Mux8~13_combout  = (instruction_D[22] & ((\Mux8~12_combout  & (\rfile[7][23]~q )) # (!\Mux8~12_combout  & ((\rfile[6][23]~q ))))) # (!instruction_D[22] & (\Mux8~12_combout ))

	.dataa(instruction_D_22),
	.datab(\Mux8~12_combout ),
	.datac(\rfile[7][23]~q ),
	.datad(\rfile[6][23]~q ),
	.cin(gnd),
	.combout(\Mux8~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~13 .lut_mask = 16'hE6C4;
defparam \Mux8~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N14
cycloneive_lcell_comb \Mux8~16 (
// Equation(s):
// \Mux8~16_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\Mux8~13_combout ))) # (!instruction_D[23] & (\Mux8~15_combout ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux8~15_combout ),
	.datad(\Mux8~13_combout ),
	.cin(gnd),
	.combout(\Mux8~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~16 .lut_mask = 16'hDC98;
defparam \Mux8~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N24
cycloneive_lcell_comb \Mux8~10 (
// Equation(s):
// \Mux8~10_combout  = (instruction_D[22] & (((\rfile[10][23]~q ) # (instruction_D[21])))) # (!instruction_D[22] & (\rfile[8][23]~q  & ((!instruction_D[21]))))

	.dataa(\rfile[8][23]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[10][23]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux8~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~10 .lut_mask = 16'hCCE2;
defparam \Mux8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N22
cycloneive_lcell_comb \Mux8~11 (
// Equation(s):
// \Mux8~11_combout  = (instruction_D[21] & ((\Mux8~10_combout  & ((\rfile[11][23]~q ))) # (!\Mux8~10_combout  & (\rfile[9][23]~q )))) # (!instruction_D[21] & (((\Mux8~10_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[9][23]~q ),
	.datac(\rfile[11][23]~q ),
	.datad(\Mux8~10_combout ),
	.cin(gnd),
	.combout(\Mux8~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~11 .lut_mask = 16'hF588;
defparam \Mux8~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N12
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[25][22]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[17][22]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[25][22]~q ),
	.datad(\rfile[17][22]~q ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hB9A8;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N26
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (instruction_D[23] & ((\Mux9~0_combout  & (\rfile[29][22]~q )) # (!\Mux9~0_combout  & ((\rfile[21][22]~q ))))) # (!instruction_D[23] & (((\Mux9~0_combout ))))

	.dataa(\rfile[29][22]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[21][22]~q ),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hBBC0;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N12
cycloneive_lcell_comb \Mux9~7 (
// Equation(s):
// \Mux9~7_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[27][22]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[19][22]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[27][22]~q ),
	.datad(\rfile[19][22]~q ),
	.cin(gnd),
	.combout(\Mux9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~7 .lut_mask = 16'hB9A8;
defparam \Mux9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N0
cycloneive_lcell_comb \Mux9~8 (
// Equation(s):
// \Mux9~8_combout  = (instruction_D[23] & ((\Mux9~7_combout  & (\rfile[31][22]~q )) # (!\Mux9~7_combout  & ((\rfile[23][22]~q ))))) # (!instruction_D[23] & (((\Mux9~7_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[31][22]~q ),
	.datac(\rfile[23][22]~q ),
	.datad(\Mux9~7_combout ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~8 .lut_mask = 16'hDDA0;
defparam \Mux9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N28
cycloneive_lcell_comb \Mux9~2 (
// Equation(s):
// \Mux9~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[22][22]~q ))) # (!instruction_D[23] & (\rfile[18][22]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][22]~q ),
	.datad(\rfile[22][22]~q ),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~2 .lut_mask = 16'hDC98;
defparam \Mux9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N24
cycloneive_lcell_comb \Mux9~3 (
// Equation(s):
// \Mux9~3_combout  = (instruction_D[24] & ((\Mux9~2_combout  & ((\rfile[30][22]~q ))) # (!\Mux9~2_combout  & (\rfile[26][22]~q )))) # (!instruction_D[24] & (((\Mux9~2_combout ))))

	.dataa(\rfile[26][22]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[30][22]~q ),
	.datad(\Mux9~2_combout ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~3 .lut_mask = 16'hF388;
defparam \Mux9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N6
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[20][22]~q )) # (!instruction_D[23] & ((\rfile[16][22]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[20][22]~q ),
	.datad(\rfile[16][22]~q ),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hD9C8;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y30_N26
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// \Mux9~5_combout  = (instruction_D[24] & ((\Mux9~4_combout  & (\rfile[28][22]~q )) # (!\Mux9~4_combout  & ((\rfile[24][22]~q ))))) # (!instruction_D[24] & (((\Mux9~4_combout ))))

	.dataa(\rfile[28][22]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[24][22]~q ),
	.datad(\Mux9~4_combout ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hBBC0;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N0
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// \Mux9~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux9~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & ((\Mux9~5_combout ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux9~3_combout ),
	.datad(\Mux9~5_combout ),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'hB9A8;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N18
cycloneive_lcell_comb \Mux9~17 (
// Equation(s):
// \Mux9~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][22]~q ))) # (!instruction_D[21] & (\rfile[12][22]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][22]~q ),
	.datad(\rfile[13][22]~q ),
	.cin(gnd),
	.combout(\Mux9~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~17 .lut_mask = 16'hDC98;
defparam \Mux9~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N18
cycloneive_lcell_comb \Mux9~18 (
// Equation(s):
// \Mux9~18_combout  = (\Mux9~17_combout  & ((\rfile[15][22]~q ) # ((!instruction_D[22])))) # (!\Mux9~17_combout  & (((instruction_D[22] & \rfile[14][22]~q ))))

	.dataa(\rfile[15][22]~q ),
	.datab(\Mux9~17_combout ),
	.datac(instruction_D_22),
	.datad(\rfile[14][22]~q ),
	.cin(gnd),
	.combout(\Mux9~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~18 .lut_mask = 16'hBC8C;
defparam \Mux9~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N24
cycloneive_lcell_comb \Mux9~10 (
// Equation(s):
// \Mux9~10_combout  = (instruction_D[21] & ((instruction_D[22]) # ((\rfile[5][22]~q )))) # (!instruction_D[21] & (!instruction_D[22] & ((\rfile[4][22]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[5][22]~q ),
	.datad(\rfile[4][22]~q ),
	.cin(gnd),
	.combout(\Mux9~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~10 .lut_mask = 16'hB9A8;
defparam \Mux9~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N10
cycloneive_lcell_comb \Mux9~11 (
// Equation(s):
// \Mux9~11_combout  = (instruction_D[22] & ((\Mux9~10_combout  & ((\rfile[7][22]~q ))) # (!\Mux9~10_combout  & (\rfile[6][22]~q )))) # (!instruction_D[22] & (((\Mux9~10_combout ))))

	.dataa(\rfile[6][22]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[7][22]~q ),
	.datad(\Mux9~10_combout ),
	.cin(gnd),
	.combout(\Mux9~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~11 .lut_mask = 16'hF388;
defparam \Mux9~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N2
cycloneive_lcell_comb \Mux9~14 (
// Equation(s):
// \Mux9~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][22]~q )) # (!instruction_D[22] & ((\rfile[1][22]~q )))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[3][22]~q ),
	.datad(\rfile[1][22]~q ),
	.cin(gnd),
	.combout(\Mux9~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~14 .lut_mask = 16'hC480;
defparam \Mux9~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N8
cycloneive_lcell_comb \Mux9~15 (
// Equation(s):
// \Mux9~15_combout  = (\Mux9~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][22]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[2][22]~q ),
	.datad(\Mux9~14_combout ),
	.cin(gnd),
	.combout(\Mux9~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~15 .lut_mask = 16'hFF20;
defparam \Mux9~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N28
cycloneive_lcell_comb \Mux9~12 (
// Equation(s):
// \Mux9~12_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][22]~q )))) # (!instruction_D[22] & (!instruction_D[21] & ((\rfile[8][22]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[10][22]~q ),
	.datad(\rfile[8][22]~q ),
	.cin(gnd),
	.combout(\Mux9~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~12 .lut_mask = 16'hB9A8;
defparam \Mux9~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N30
cycloneive_lcell_comb \Mux9~13 (
// Equation(s):
// \Mux9~13_combout  = (instruction_D[21] & ((\Mux9~12_combout  & (\rfile[11][22]~q )) # (!\Mux9~12_combout  & ((\rfile[9][22]~q ))))) # (!instruction_D[21] & (((\Mux9~12_combout ))))

	.dataa(instruction_D_21),
	.datab(\rfile[11][22]~q ),
	.datac(\rfile[9][22]~q ),
	.datad(\Mux9~12_combout ),
	.cin(gnd),
	.combout(\Mux9~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~13 .lut_mask = 16'hDDA0;
defparam \Mux9~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N12
cycloneive_lcell_comb \Mux9~16 (
// Equation(s):
// \Mux9~16_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\Mux9~13_combout ))) # (!instruction_D[24] & (\Mux9~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux9~15_combout ),
	.datad(\Mux9~13_combout ),
	.cin(gnd),
	.combout(\Mux9~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~16 .lut_mask = 16'hDC98;
defparam \Mux9~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N28
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[21][21]~q ))) # (!instruction_D[23] & (\rfile[17][21]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[17][21]~q ),
	.datad(\rfile[21][21]~q ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hDC98;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N8
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (instruction_D[24] & ((\Mux10~0_combout  & ((\rfile[29][21]~q ))) # (!\Mux10~0_combout  & (\rfile[25][21]~q )))) # (!instruction_D[24] & (((\Mux10~0_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[25][21]~q ),
	.datac(\rfile[29][21]~q ),
	.datad(\Mux10~0_combout ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hF588;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N28
cycloneive_lcell_comb \Mux10~7 (
// Equation(s):
// \Mux10~7_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[23][21]~q )) # (!instruction_D[23] & ((\rfile[19][21]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[23][21]~q ),
	.datad(\rfile[19][21]~q ),
	.cin(gnd),
	.combout(\Mux10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~7 .lut_mask = 16'hD9C8;
defparam \Mux10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N8
cycloneive_lcell_comb \Mux10~8 (
// Equation(s):
// \Mux10~8_combout  = (\Mux10~7_combout  & ((\rfile[31][21]~q ) # ((!instruction_D[24])))) # (!\Mux10~7_combout  & (((\rfile[27][21]~q  & instruction_D[24]))))

	.dataa(\rfile[31][21]~q ),
	.datab(\Mux10~7_combout ),
	.datac(\rfile[27][21]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~8 .lut_mask = 16'hB8CC;
defparam \Mux10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y33_N27
dffeas \rfile[20][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][21] .is_wysiwyg = "true";
defparam \rfile[20][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N6
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\rfile[24][21]~q ))) # (!instruction_D[24] & (\rfile[16][21]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[16][21]~q ),
	.datad(\rfile[24][21]~q ),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hDC98;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N26
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// \Mux10~5_combout  = (instruction_D[23] & ((\Mux10~4_combout  & (\rfile[28][21]~q )) # (!\Mux10~4_combout  & ((\rfile[20][21]~q ))))) # (!instruction_D[23] & (((\Mux10~4_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[28][21]~q ),
	.datac(\rfile[20][21]~q ),
	.datad(\Mux10~4_combout ),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hDDA0;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N24
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][21]~q )))) # (!instruction_D[24] & (!instruction_D[23] & ((\rfile[18][21]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[26][21]~q ),
	.datad(\rfile[18][21]~q ),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hB9A8;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N2
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (instruction_D[23] & ((\Mux10~2_combout  & ((\rfile[30][21]~q ))) # (!\Mux10~2_combout  & (\rfile[22][21]~q )))) # (!instruction_D[23] & (((\Mux10~2_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[22][21]~q ),
	.datac(\rfile[30][21]~q ),
	.datad(\Mux10~2_combout ),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'hF588;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N0
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// \Mux10~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux10~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & (\Mux10~5_combout )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux10~5_combout ),
	.datad(\Mux10~3_combout ),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'hBA98;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N1
dffeas \rfile[4][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][21] .is_wysiwyg = "true";
defparam \rfile[4][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N0
cycloneive_lcell_comb \Mux10~12 (
// Equation(s):
// \Mux10~12_combout  = (instruction_D[21] & ((\rfile[5][21]~q ) # ((instruction_D[22])))) # (!instruction_D[21] & (((\rfile[4][21]~q  & !instruction_D[22]))))

	.dataa(instruction_D_21),
	.datab(\rfile[5][21]~q ),
	.datac(\rfile[4][21]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux10~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~12 .lut_mask = 16'hAAD8;
defparam \Mux10~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N26
cycloneive_lcell_comb \Mux10~13 (
// Equation(s):
// \Mux10~13_combout  = (instruction_D[22] & ((\Mux10~12_combout  & ((\rfile[7][21]~q ))) # (!\Mux10~12_combout  & (\rfile[6][21]~q )))) # (!instruction_D[22] & (((\Mux10~12_combout ))))

	.dataa(\rfile[6][21]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[7][21]~q ),
	.datad(\Mux10~12_combout ),
	.cin(gnd),
	.combout(\Mux10~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~13 .lut_mask = 16'hF388;
defparam \Mux10~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N10
cycloneive_lcell_comb \Mux10~14 (
// Equation(s):
// \Mux10~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][21]~q ))) # (!instruction_D[22] & (\rfile[1][21]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[1][21]~q ),
	.datad(\rfile[3][21]~q ),
	.cin(gnd),
	.combout(\Mux10~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~14 .lut_mask = 16'hA820;
defparam \Mux10~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N10
cycloneive_lcell_comb \Mux10~15 (
// Equation(s):
// \Mux10~15_combout  = (\Mux10~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][21]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[2][21]~q ),
	.datad(\Mux10~14_combout ),
	.cin(gnd),
	.combout(\Mux10~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~15 .lut_mask = 16'hFF20;
defparam \Mux10~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N30
cycloneive_lcell_comb \Mux10~16 (
// Equation(s):
// \Mux10~16_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\Mux10~13_combout )) # (!instruction_D[23] & ((\Mux10~15_combout )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux10~13_combout ),
	.datad(\Mux10~15_combout ),
	.cin(gnd),
	.combout(\Mux10~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~16 .lut_mask = 16'hD9C8;
defparam \Mux10~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N30
cycloneive_lcell_comb \Mux10~17 (
// Equation(s):
// \Mux10~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][21]~q ))) # (!instruction_D[21] & (\rfile[12][21]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][21]~q ),
	.datad(\rfile[13][21]~q ),
	.cin(gnd),
	.combout(\Mux10~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~17 .lut_mask = 16'hDC98;
defparam \Mux10~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N16
cycloneive_lcell_comb \Mux10~18 (
// Equation(s):
// \Mux10~18_combout  = (instruction_D[22] & ((\Mux10~17_combout  & ((\rfile[15][21]~q ))) # (!\Mux10~17_combout  & (\rfile[14][21]~q )))) # (!instruction_D[22] & (((\Mux10~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[14][21]~q ),
	.datac(\Mux10~17_combout ),
	.datad(\rfile[15][21]~q ),
	.cin(gnd),
	.combout(\Mux10~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~18 .lut_mask = 16'hF858;
defparam \Mux10~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N0
cycloneive_lcell_comb \Mux10~10 (
// Equation(s):
// \Mux10~10_combout  = (instruction_D[21] & (((instruction_D[22])))) # (!instruction_D[21] & ((instruction_D[22] & ((\rfile[10][21]~q ))) # (!instruction_D[22] & (\rfile[8][21]~q ))))

	.dataa(\rfile[8][21]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[10][21]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux10~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~10 .lut_mask = 16'hFC22;
defparam \Mux10~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N24
cycloneive_lcell_comb \Mux10~11 (
// Equation(s):
// \Mux10~11_combout  = (instruction_D[21] & ((\Mux10~10_combout  & ((\rfile[11][21]~q ))) # (!\Mux10~10_combout  & (\rfile[9][21]~q )))) # (!instruction_D[21] & (((\Mux10~10_combout ))))

	.dataa(\rfile[9][21]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[11][21]~q ),
	.datad(\Mux10~10_combout ),
	.cin(gnd),
	.combout(\Mux10~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~11 .lut_mask = 16'hF388;
defparam \Mux10~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y29_N28
cycloneive_lcell_comb \Mux11~7 (
// Equation(s):
// \Mux11~7_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[27][20]~q )) # (!instruction_D[24] & ((\rfile[19][20]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[27][20]~q ),
	.datad(\rfile[19][20]~q ),
	.cin(gnd),
	.combout(\Mux11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~7 .lut_mask = 16'hD9C8;
defparam \Mux11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N20
cycloneive_lcell_comb \Mux11~8 (
// Equation(s):
// \Mux11~8_combout  = (instruction_D[23] & ((\Mux11~7_combout  & (\rfile[31][20]~q )) # (!\Mux11~7_combout  & ((\rfile[23][20]~q ))))) # (!instruction_D[23] & (((\Mux11~7_combout ))))

	.dataa(\rfile[31][20]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[23][20]~q ),
	.datad(\Mux11~7_combout ),
	.cin(gnd),
	.combout(\Mux11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~8 .lut_mask = 16'hBBC0;
defparam \Mux11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y35_N27
dffeas \rfile[22][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][20] .is_wysiwyg = "true";
defparam \rfile[22][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N26
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[22][20]~q )) # (!instruction_D[23] & ((\rfile[18][20]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[22][20]~q ),
	.datad(\rfile[18][20]~q ),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hD9C8;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N16
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (instruction_D[24] & ((\Mux11~2_combout  & ((\rfile[30][20]~q ))) # (!\Mux11~2_combout  & (\rfile[26][20]~q )))) # (!instruction_D[24] & (((\Mux11~2_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[26][20]~q ),
	.datac(\rfile[30][20]~q ),
	.datad(\Mux11~2_combout ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hF588;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y33_N5
dffeas \rfile[24][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[24][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[24][20] .is_wysiwyg = "true";
defparam \rfile[24][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X76_Y33_N18
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[20][20]~q ))) # (!instruction_D[23] & (\rfile[16][20]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[16][20]~q ),
	.datad(\rfile[20][20]~q ),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hDC98;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N4
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// \Mux11~5_combout  = (instruction_D[24] & ((\Mux11~4_combout  & (\rfile[28][20]~q )) # (!\Mux11~4_combout  & ((\rfile[24][20]~q ))))) # (!instruction_D[24] & (((\Mux11~4_combout ))))

	.dataa(\rfile[28][20]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[24][20]~q ),
	.datad(\Mux11~4_combout ),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hBBC0;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N22
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// \Mux11~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\Mux11~3_combout )) # (!instruction_D[22] & ((\Mux11~5_combout )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux11~3_combout ),
	.datad(\Mux11~5_combout ),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'hD9C8;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y28_N27
dffeas \rfile[25][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[25][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[25][20] .is_wysiwyg = "true";
defparam \rfile[25][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N26
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (instruction_D[24] & (((\rfile[25][20]~q ) # (instruction_D[23])))) # (!instruction_D[24] & (\rfile[17][20]~q  & ((!instruction_D[23]))))

	.dataa(instruction_D_24),
	.datab(\rfile[17][20]~q ),
	.datac(\rfile[25][20]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hAAE4;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N26
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (instruction_D[23] & ((\Mux11~0_combout  & (\rfile[29][20]~q )) # (!\Mux11~0_combout  & ((\rfile[21][20]~q ))))) # (!instruction_D[23] & (\Mux11~0_combout ))

	.dataa(instruction_D_23),
	.datab(\Mux11~0_combout ),
	.datac(\rfile[29][20]~q ),
	.datad(\rfile[21][20]~q ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hE6C4;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N19
dffeas \rfile[1][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[1][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[1][20] .is_wysiwyg = "true";
defparam \rfile[1][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N18
cycloneive_lcell_comb \Mux11~14 (
// Equation(s):
// \Mux11~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][20]~q ))) # (!instruction_D[22] & (\rfile[1][20]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[1][20]~q ),
	.datad(\rfile[3][20]~q ),
	.cin(gnd),
	.combout(\Mux11~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~14 .lut_mask = 16'hA820;
defparam \Mux11~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N26
cycloneive_lcell_comb \Mux11~15 (
// Equation(s):
// \Mux11~15_combout  = (\Mux11~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][20]~q )))

	.dataa(instruction_D_22),
	.datab(\Mux11~14_combout ),
	.datac(instruction_D_21),
	.datad(\rfile[2][20]~q ),
	.cin(gnd),
	.combout(\Mux11~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~15 .lut_mask = 16'hCECC;
defparam \Mux11~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N16
cycloneive_lcell_comb \Mux11~12 (
// Equation(s):
// \Mux11~12_combout  = (instruction_D[22] & (((\rfile[10][20]~q ) # (instruction_D[21])))) # (!instruction_D[22] & (\rfile[8][20]~q  & ((!instruction_D[21]))))

	.dataa(\rfile[8][20]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[10][20]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux11~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~12 .lut_mask = 16'hCCE2;
defparam \Mux11~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N5
dffeas \rfile[11][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[11][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[11][20] .is_wysiwyg = "true";
defparam \rfile[11][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N4
cycloneive_lcell_comb \Mux11~13 (
// Equation(s):
// \Mux11~13_combout  = (instruction_D[21] & ((\Mux11~12_combout  & (\rfile[11][20]~q )) # (!\Mux11~12_combout  & ((\rfile[9][20]~q ))))) # (!instruction_D[21] & (\Mux11~12_combout ))

	.dataa(instruction_D_21),
	.datab(\Mux11~12_combout ),
	.datac(\rfile[11][20]~q ),
	.datad(\rfile[9][20]~q ),
	.cin(gnd),
	.combout(\Mux11~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~13 .lut_mask = 16'hE6C4;
defparam \Mux11~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N8
cycloneive_lcell_comb \Mux11~16 (
// Equation(s):
// \Mux11~16_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\Mux11~13_combout ))) # (!instruction_D[24] & (\Mux11~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux11~15_combout ),
	.datad(\Mux11~13_combout ),
	.cin(gnd),
	.combout(\Mux11~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~16 .lut_mask = 16'hDC98;
defparam \Mux11~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N14
cycloneive_lcell_comb \Mux11~17 (
// Equation(s):
// \Mux11~17_combout  = (instruction_D[21] & ((\rfile[13][20]~q ) # ((instruction_D[22])))) # (!instruction_D[21] & (((!instruction_D[22] & \rfile[12][20]~q ))))

	.dataa(instruction_D_21),
	.datab(\rfile[13][20]~q ),
	.datac(instruction_D_22),
	.datad(\rfile[12][20]~q ),
	.cin(gnd),
	.combout(\Mux11~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~17 .lut_mask = 16'hADA8;
defparam \Mux11~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N18
cycloneive_lcell_comb \Mux11~18 (
// Equation(s):
// \Mux11~18_combout  = (instruction_D[22] & ((\Mux11~17_combout  & (\rfile[15][20]~q )) # (!\Mux11~17_combout  & ((\rfile[14][20]~q ))))) # (!instruction_D[22] & (((\Mux11~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[15][20]~q ),
	.datac(\rfile[14][20]~q ),
	.datad(\Mux11~17_combout ),
	.cin(gnd),
	.combout(\Mux11~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~18 .lut_mask = 16'hDDA0;
defparam \Mux11~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N10
cycloneive_lcell_comb \Mux11~10 (
// Equation(s):
// \Mux11~10_combout  = (instruction_D[21] & ((instruction_D[22]) # ((\rfile[5][20]~q )))) # (!instruction_D[21] & (!instruction_D[22] & ((\rfile[4][20]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[5][20]~q ),
	.datad(\rfile[4][20]~q ),
	.cin(gnd),
	.combout(\Mux11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~10 .lut_mask = 16'hB9A8;
defparam \Mux11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N6
cycloneive_lcell_comb \Mux11~11 (
// Equation(s):
// \Mux11~11_combout  = (instruction_D[22] & ((\Mux11~10_combout  & ((\rfile[7][20]~q ))) # (!\Mux11~10_combout  & (\rfile[6][20]~q )))) # (!instruction_D[22] & (((\Mux11~10_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[6][20]~q ),
	.datac(\rfile[7][20]~q ),
	.datad(\Mux11~10_combout ),
	.cin(gnd),
	.combout(\Mux11~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~11 .lut_mask = 16'hF588;
defparam \Mux11~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y29_N12
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// \Mux12~7_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[23][19]~q ))) # (!instruction_D[23] & (\rfile[19][19]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[19][19]~q ),
	.datad(\rfile[23][19]~q ),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hDC98;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N10
cycloneive_lcell_comb \Mux12~8 (
// Equation(s):
// \Mux12~8_combout  = (instruction_D[24] & ((\Mux12~7_combout  & ((\rfile[31][19]~q ))) # (!\Mux12~7_combout  & (\rfile[27][19]~q )))) # (!instruction_D[24] & (\Mux12~7_combout ))

	.dataa(instruction_D_24),
	.datab(\Mux12~7_combout ),
	.datac(\rfile[27][19]~q ),
	.datad(\rfile[31][19]~q ),
	.cin(gnd),
	.combout(\Mux12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~8 .lut_mask = 16'hEC64;
defparam \Mux12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N22
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[21][19]~q ))) # (!instruction_D[23] & (\rfile[17][19]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[17][19]~q ),
	.datad(\rfile[21][19]~q ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hDC98;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N12
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (instruction_D[24] & ((\Mux12~0_combout  & ((\rfile[29][19]~q ))) # (!\Mux12~0_combout  & (\rfile[25][19]~q )))) # (!instruction_D[24] & (((\Mux12~0_combout ))))

	.dataa(\rfile[25][19]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[29][19]~q ),
	.datad(\Mux12~0_combout ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hF388;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N6
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[26][19]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[18][19]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][19]~q ),
	.datad(\rfile[26][19]~q ),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'hBA98;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N14
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// \Mux12~3_combout  = (instruction_D[23] & ((\Mux12~2_combout  & ((\rfile[30][19]~q ))) # (!\Mux12~2_combout  & (\rfile[22][19]~q )))) # (!instruction_D[23] & (((\Mux12~2_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[22][19]~q ),
	.datac(\rfile[30][19]~q ),
	.datad(\Mux12~2_combout ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'hF588;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N2
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[24][19]~q )) # (!instruction_D[24] & ((\rfile[16][19]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[24][19]~q ),
	.datad(\rfile[16][19]~q ),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'hD9C8;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N28
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// \Mux12~5_combout  = (instruction_D[23] & ((\Mux12~4_combout  & (\rfile[28][19]~q )) # (!\Mux12~4_combout  & ((\rfile[20][19]~q ))))) # (!instruction_D[23] & (((\Mux12~4_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[28][19]~q ),
	.datac(\rfile[20][19]~q ),
	.datad(\Mux12~4_combout ),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hDDA0;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N18
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// \Mux12~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & (\Mux12~3_combout )) # (!instruction_D[22] & ((\Mux12~5_combout )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux12~3_combout ),
	.datad(\Mux12~5_combout ),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'hD9C8;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N10
cycloneive_lcell_comb \Mux12~17 (
// Equation(s):
// \Mux12~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][19]~q ))) # (!instruction_D[21] & (\rfile[12][19]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][19]~q ),
	.datad(\rfile[13][19]~q ),
	.cin(gnd),
	.combout(\Mux12~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~17 .lut_mask = 16'hDC98;
defparam \Mux12~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N2
cycloneive_lcell_comb \Mux12~18 (
// Equation(s):
// \Mux12~18_combout  = (instruction_D[22] & ((\Mux12~17_combout  & ((\rfile[15][19]~q ))) # (!\Mux12~17_combout  & (\rfile[14][19]~q )))) # (!instruction_D[22] & (((\Mux12~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[14][19]~q ),
	.datac(\rfile[15][19]~q ),
	.datad(\Mux12~17_combout ),
	.cin(gnd),
	.combout(\Mux12~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~18 .lut_mask = 16'hF588;
defparam \Mux12~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N12
cycloneive_lcell_comb \Mux12~10 (
// Equation(s):
// \Mux12~10_combout  = (instruction_D[21] & (((instruction_D[22])))) # (!instruction_D[21] & ((instruction_D[22] & ((\rfile[10][19]~q ))) # (!instruction_D[22] & (\rfile[8][19]~q ))))

	.dataa(\rfile[8][19]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[10][19]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux12~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~10 .lut_mask = 16'hFC22;
defparam \Mux12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N18
cycloneive_lcell_comb \Mux12~11 (
// Equation(s):
// \Mux12~11_combout  = (instruction_D[21] & ((\Mux12~10_combout  & ((\rfile[11][19]~q ))) # (!\Mux12~10_combout  & (\rfile[9][19]~q )))) # (!instruction_D[21] & (\Mux12~10_combout ))

	.dataa(instruction_D_21),
	.datab(\Mux12~10_combout ),
	.datac(\rfile[9][19]~q ),
	.datad(\rfile[11][19]~q ),
	.cin(gnd),
	.combout(\Mux12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~11 .lut_mask = 16'hEC64;
defparam \Mux12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N21
dffeas \rfile[4][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[4][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[4][19] .is_wysiwyg = "true";
defparam \rfile[4][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N3
dffeas \rfile[5][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[5][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[5][19] .is_wysiwyg = "true";
defparam \rfile[5][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N20
cycloneive_lcell_comb \Mux12~12 (
// Equation(s):
// \Mux12~12_combout  = (instruction_D[21] & ((instruction_D[22]) # ((\rfile[5][19]~q )))) # (!instruction_D[21] & (!instruction_D[22] & (\rfile[4][19]~q )))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[4][19]~q ),
	.datad(\rfile[5][19]~q ),
	.cin(gnd),
	.combout(\Mux12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~12 .lut_mask = 16'hBA98;
defparam \Mux12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N2
cycloneive_lcell_comb \Mux12~13 (
// Equation(s):
// \Mux12~13_combout  = (instruction_D[22] & ((\Mux12~12_combout  & ((\rfile[7][19]~q ))) # (!\Mux12~12_combout  & (\rfile[6][19]~q )))) # (!instruction_D[22] & (((\Mux12~12_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[6][19]~q ),
	.datac(\rfile[7][19]~q ),
	.datad(\Mux12~12_combout ),
	.cin(gnd),
	.combout(\Mux12~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~13 .lut_mask = 16'hF588;
defparam \Mux12~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N24
cycloneive_lcell_comb \Mux12~14 (
// Equation(s):
// \Mux12~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][19]~q )) # (!instruction_D[22] & ((\rfile[1][19]~q )))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[3][19]~q ),
	.datad(\rfile[1][19]~q ),
	.cin(gnd),
	.combout(\Mux12~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~14 .lut_mask = 16'hA280;
defparam \Mux12~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N2
cycloneive_lcell_comb \Mux12~15 (
// Equation(s):
// \Mux12~15_combout  = (\Mux12~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][19]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[2][19]~q ),
	.datad(\Mux12~14_combout ),
	.cin(gnd),
	.combout(\Mux12~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~15 .lut_mask = 16'hFF20;
defparam \Mux12~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N10
cycloneive_lcell_comb \Mux12~16 (
// Equation(s):
// \Mux12~16_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\Mux12~13_combout )))) # (!instruction_D[23] & (!instruction_D[24] & ((\Mux12~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux12~13_combout ),
	.datad(\Mux12~15_combout ),
	.cin(gnd),
	.combout(\Mux12~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~16 .lut_mask = 16'hB9A8;
defparam \Mux12~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y28_N18
cycloneive_lcell_comb \Mux13~7 (
// Equation(s):
// \Mux13~7_combout  = (instruction_D[24] & (((instruction_D[23]) # (\rfile[27][18]~q )))) # (!instruction_D[24] & (\rfile[19][18]~q  & (!instruction_D[23])))

	.dataa(instruction_D_24),
	.datab(\rfile[19][18]~q ),
	.datac(instruction_D_23),
	.datad(\rfile[27][18]~q ),
	.cin(gnd),
	.combout(\Mux13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~7 .lut_mask = 16'hAEA4;
defparam \Mux13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N30
cycloneive_lcell_comb \Mux13~8 (
// Equation(s):
// \Mux13~8_combout  = (instruction_D[23] & ((\Mux13~7_combout  & ((\rfile[31][18]~q ))) # (!\Mux13~7_combout  & (\rfile[23][18]~q )))) # (!instruction_D[23] & (((\Mux13~7_combout ))))

	.dataa(\rfile[23][18]~q ),
	.datab(instruction_D_23),
	.datac(\Mux13~7_combout ),
	.datad(\rfile[31][18]~q ),
	.cin(gnd),
	.combout(\Mux13~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~8 .lut_mask = 16'hF838;
defparam \Mux13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N12
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & (\rfile[25][18]~q )) # (!instruction_D[24] & ((\rfile[17][18]~q )))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[25][18]~q ),
	.datad(\rfile[17][18]~q ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hD9C8;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N14
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (instruction_D[23] & ((\Mux13~0_combout  & ((\rfile[29][18]~q ))) # (!\Mux13~0_combout  & (\rfile[21][18]~q )))) # (!instruction_D[23] & (((\Mux13~0_combout ))))

	.dataa(\rfile[21][18]~q ),
	.datab(\rfile[29][18]~q ),
	.datac(instruction_D_23),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hCFA0;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y35_N22
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & ((\rfile[22][18]~q ))) # (!instruction_D[23] & (\rfile[18][18]~q ))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[18][18]~q ),
	.datad(\rfile[22][18]~q ),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'hDC98;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N4
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (instruction_D[24] & ((\Mux13~2_combout  & ((\rfile[30][18]~q ))) # (!\Mux13~2_combout  & (\rfile[26][18]~q )))) # (!instruction_D[24] & (((\Mux13~2_combout ))))

	.dataa(\rfile[26][18]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[30][18]~q ),
	.datad(\Mux13~2_combout ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'hF388;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N12
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[20][18]~q )) # (!instruction_D[23] & ((\rfile[16][18]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[20][18]~q ),
	.datad(\rfile[16][18]~q ),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hD9C8;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y33_N10
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// \Mux13~5_combout  = (instruction_D[24] & ((\Mux13~4_combout  & ((\rfile[28][18]~q ))) # (!\Mux13~4_combout  & (\rfile[24][18]~q )))) # (!instruction_D[24] & (((\Mux13~4_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[24][18]~q ),
	.datac(\rfile[28][18]~q ),
	.datad(\Mux13~4_combout ),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hF588;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N24
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// \Mux13~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux13~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & ((\Mux13~5_combout ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux13~3_combout ),
	.datad(\Mux13~5_combout ),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'hB9A8;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N4
cycloneive_lcell_comb \Mux13~10 (
// Equation(s):
// \Mux13~10_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & (\rfile[5][18]~q )) # (!instruction_D[21] & ((\rfile[4][18]~q )))))

	.dataa(\rfile[5][18]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[4][18]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux13~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~10 .lut_mask = 16'hEE30;
defparam \Mux13~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N20
cycloneive_lcell_comb \Mux13~11 (
// Equation(s):
// \Mux13~11_combout  = (instruction_D[22] & ((\Mux13~10_combout  & ((\rfile[7][18]~q ))) # (!\Mux13~10_combout  & (\rfile[6][18]~q )))) # (!instruction_D[22] & (((\Mux13~10_combout ))))

	.dataa(\rfile[6][18]~q ),
	.datab(\rfile[7][18]~q ),
	.datac(instruction_D_22),
	.datad(\Mux13~10_combout ),
	.cin(gnd),
	.combout(\Mux13~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~11 .lut_mask = 16'hCFA0;
defparam \Mux13~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N6
cycloneive_lcell_comb \Mux13~17 (
// Equation(s):
// \Mux13~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][18]~q ))) # (!instruction_D[21] & (\rfile[12][18]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][18]~q ),
	.datad(\rfile[13][18]~q ),
	.cin(gnd),
	.combout(\Mux13~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~17 .lut_mask = 16'hDC98;
defparam \Mux13~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N4
cycloneive_lcell_comb \Mux13~18 (
// Equation(s):
// \Mux13~18_combout  = (instruction_D[22] & ((\Mux13~17_combout  & ((\rfile[15][18]~q ))) # (!\Mux13~17_combout  & (\rfile[14][18]~q )))) # (!instruction_D[22] & (((\Mux13~17_combout ))))

	.dataa(\rfile[14][18]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[15][18]~q ),
	.datad(\Mux13~17_combout ),
	.cin(gnd),
	.combout(\Mux13~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~18 .lut_mask = 16'hF388;
defparam \Mux13~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N14
cycloneive_lcell_comb \Mux13~14 (
// Equation(s):
// \Mux13~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][18]~q ))) # (!instruction_D[22] & (\rfile[1][18]~q ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[1][18]~q ),
	.datad(\rfile[3][18]~q ),
	.cin(gnd),
	.combout(\Mux13~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~14 .lut_mask = 16'hA820;
defparam \Mux13~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N26
cycloneive_lcell_comb \Mux13~15 (
// Equation(s):
// \Mux13~15_combout  = (\Mux13~14_combout ) # ((instruction_D[22] & (!instruction_D[21] & \rfile[2][18]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux13~14_combout ),
	.datad(\rfile[2][18]~q ),
	.cin(gnd),
	.combout(\Mux13~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~15 .lut_mask = 16'hF2F0;
defparam \Mux13~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N16
cycloneive_lcell_comb \Mux13~12 (
// Equation(s):
// \Mux13~12_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][18]~q )))) # (!instruction_D[22] & (!instruction_D[21] & (\rfile[8][18]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[8][18]~q ),
	.datad(\rfile[10][18]~q ),
	.cin(gnd),
	.combout(\Mux13~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~12 .lut_mask = 16'hBA98;
defparam \Mux13~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N18
cycloneive_lcell_comb \Mux13~13 (
// Equation(s):
// \Mux13~13_combout  = (instruction_D[21] & ((\Mux13~12_combout  & ((\rfile[11][18]~q ))) # (!\Mux13~12_combout  & (\rfile[9][18]~q )))) # (!instruction_D[21] & (((\Mux13~12_combout ))))

	.dataa(\rfile[9][18]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[11][18]~q ),
	.datad(\Mux13~12_combout ),
	.cin(gnd),
	.combout(\Mux13~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~13 .lut_mask = 16'hF388;
defparam \Mux13~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N16
cycloneive_lcell_comb \Mux13~16 (
// Equation(s):
// \Mux13~16_combout  = (instruction_D[23] & (instruction_D[24])) # (!instruction_D[23] & ((instruction_D[24] & ((\Mux13~13_combout ))) # (!instruction_D[24] & (\Mux13~15_combout ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\Mux13~15_combout ),
	.datad(\Mux13~13_combout ),
	.cin(gnd),
	.combout(\Mux13~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~16 .lut_mask = 16'hDC98;
defparam \Mux13~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N6
cycloneive_lcell_comb \rfile[20][17]~feeder (
// Equation(s):
// \rfile[20][17]~feeder_combout  = \wdat_WB[17]~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat_WB_17),
	.datad(gnd),
	.cin(gnd),
	.combout(\rfile[20][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \rfile[20][17]~feeder .lut_mask = 16'hF0F0;
defparam \rfile[20][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N7
dffeas \rfile[20][17] (
	.clk(!CLK),
	.d(\rfile[20][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[20][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[20][17] .is_wysiwyg = "true";
defparam \rfile[20][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y33_N0
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// \Mux14~4_combout  = (instruction_D[24] & ((\rfile[24][17]~q ) # ((instruction_D[23])))) # (!instruction_D[24] & (((\rfile[16][17]~q  & !instruction_D[23]))))

	.dataa(instruction_D_24),
	.datab(\rfile[24][17]~q ),
	.datac(\rfile[16][17]~q ),
	.datad(instruction_D_23),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hAAD8;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N14
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (instruction_D[23] & ((\Mux14~4_combout  & ((\rfile[28][17]~q ))) # (!\Mux14~4_combout  & (\rfile[20][17]~q )))) # (!instruction_D[23] & (((\Mux14~4_combout ))))

	.dataa(instruction_D_23),
	.datab(\rfile[20][17]~q ),
	.datac(\rfile[28][17]~q ),
	.datad(\Mux14~4_combout ),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hF588;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X74_Y35_N31
dffeas \rfile[22][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[22][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[22][17] .is_wysiwyg = "true";
defparam \rfile[22][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X74_Y35_N30
cycloneive_lcell_comb \Mux14~3 (
// Equation(s):
// \Mux14~3_combout  = (\Mux14~2_combout  & (((\rfile[30][17]~q )) # (!instruction_D[23]))) # (!\Mux14~2_combout  & (instruction_D[23] & (\rfile[22][17]~q )))

	.dataa(\Mux14~2_combout ),
	.datab(instruction_D_23),
	.datac(\rfile[22][17]~q ),
	.datad(\rfile[30][17]~q ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~3 .lut_mask = 16'hEA62;
defparam \Mux14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N24
cycloneive_lcell_comb \Mux14~6 (
// Equation(s):
// \Mux14~6_combout  = (instruction_D[21] & (instruction_D[22])) # (!instruction_D[21] & ((instruction_D[22] & ((\Mux14~3_combout ))) # (!instruction_D[22] & (\Mux14~5_combout ))))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\Mux14~5_combout ),
	.datad(\Mux14~3_combout ),
	.cin(gnd),
	.combout(\Mux14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~6 .lut_mask = 16'hDC98;
defparam \Mux14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y28_N28
cycloneive_lcell_comb \Mux14~7 (
// Equation(s):
// \Mux14~7_combout  = (instruction_D[23] & (((instruction_D[24]) # (\rfile[23][17]~q )))) # (!instruction_D[23] & (\rfile[19][17]~q  & (!instruction_D[24])))

	.dataa(instruction_D_23),
	.datab(\rfile[19][17]~q ),
	.datac(instruction_D_24),
	.datad(\rfile[23][17]~q ),
	.cin(gnd),
	.combout(\Mux14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~7 .lut_mask = 16'hAEA4;
defparam \Mux14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y28_N2
cycloneive_lcell_comb \Mux14~8 (
// Equation(s):
// \Mux14~8_combout  = (instruction_D[24] & ((\Mux14~7_combout  & (\rfile[31][17]~q )) # (!\Mux14~7_combout  & ((\rfile[27][17]~q ))))) # (!instruction_D[24] & (((\Mux14~7_combout ))))

	.dataa(\rfile[31][17]~q ),
	.datab(\rfile[27][17]~q ),
	.datac(instruction_D_24),
	.datad(\Mux14~7_combout ),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~8 .lut_mask = 16'hAFC0;
defparam \Mux14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N6
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (instruction_D[23] & ((instruction_D[24]) # ((\rfile[21][17]~q )))) # (!instruction_D[23] & (!instruction_D[24] & ((\rfile[17][17]~q ))))

	.dataa(instruction_D_23),
	.datab(instruction_D_24),
	.datac(\rfile[21][17]~q ),
	.datad(\rfile[17][17]~q ),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hB9A8;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N24
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (instruction_D[24] & ((\Mux14~0_combout  & ((\rfile[29][17]~q ))) # (!\Mux14~0_combout  & (\rfile[25][17]~q )))) # (!instruction_D[24] & (((\Mux14~0_combout ))))

	.dataa(\rfile[25][17]~q ),
	.datab(instruction_D_24),
	.datac(\rfile[29][17]~q ),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hF388;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N2
cycloneive_lcell_comb \Mux14~10 (
// Equation(s):
// \Mux14~10_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][17]~q )))) # (!instruction_D[22] & (!instruction_D[21] & (\rfile[8][17]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[8][17]~q ),
	.datad(\rfile[10][17]~q ),
	.cin(gnd),
	.combout(\Mux14~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~10 .lut_mask = 16'hBA98;
defparam \Mux14~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N0
cycloneive_lcell_comb \Mux14~11 (
// Equation(s):
// \Mux14~11_combout  = (instruction_D[21] & ((\Mux14~10_combout  & (\rfile[11][17]~q )) # (!\Mux14~10_combout  & ((\rfile[9][17]~q ))))) # (!instruction_D[21] & (((\Mux14~10_combout ))))

	.dataa(\rfile[11][17]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[9][17]~q ),
	.datad(\Mux14~10_combout ),
	.cin(gnd),
	.combout(\Mux14~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~11 .lut_mask = 16'hBBC0;
defparam \Mux14~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N4
cycloneive_lcell_comb \Mux14~12 (
// Equation(s):
// \Mux14~12_combout  = (instruction_D[22] & (((instruction_D[21])))) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[5][17]~q ))) # (!instruction_D[21] & (\rfile[4][17]~q ))))

	.dataa(\rfile[4][17]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[5][17]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux14~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~12 .lut_mask = 16'hFC22;
defparam \Mux14~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N28
cycloneive_lcell_comb \Mux14~13 (
// Equation(s):
// \Mux14~13_combout  = (instruction_D[22] & ((\Mux14~12_combout  & (\rfile[7][17]~q )) # (!\Mux14~12_combout  & ((\rfile[6][17]~q ))))) # (!instruction_D[22] & (\Mux14~12_combout ))

	.dataa(instruction_D_22),
	.datab(\Mux14~12_combout ),
	.datac(\rfile[7][17]~q ),
	.datad(\rfile[6][17]~q ),
	.cin(gnd),
	.combout(\Mux14~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~13 .lut_mask = 16'hE6C4;
defparam \Mux14~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N28
cycloneive_lcell_comb \Mux14~14 (
// Equation(s):
// \Mux14~14_combout  = (instruction_D[21] & ((instruction_D[22] & (\rfile[3][17]~q )) # (!instruction_D[22] & ((\rfile[1][17]~q )))))

	.dataa(\rfile[3][17]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[1][17]~q ),
	.datad(instruction_D_21),
	.cin(gnd),
	.combout(\Mux14~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~14 .lut_mask = 16'hB800;
defparam \Mux14~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N16
cycloneive_lcell_comb \Mux14~15 (
// Equation(s):
// \Mux14~15_combout  = (\Mux14~14_combout ) # ((!instruction_D[21] & (\rfile[2][17]~q  & instruction_D[22])))

	.dataa(instruction_D_21),
	.datab(\rfile[2][17]~q ),
	.datac(instruction_D_22),
	.datad(\Mux14~14_combout ),
	.cin(gnd),
	.combout(\Mux14~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~15 .lut_mask = 16'hFF40;
defparam \Mux14~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N26
cycloneive_lcell_comb \Mux14~16 (
// Equation(s):
// \Mux14~16_combout  = (instruction_D[23] & ((\Mux14~13_combout ) # ((instruction_D[24])))) # (!instruction_D[23] & (((!instruction_D[24] & \Mux14~15_combout ))))

	.dataa(instruction_D_23),
	.datab(\Mux14~13_combout ),
	.datac(instruction_D_24),
	.datad(\Mux14~15_combout ),
	.cin(gnd),
	.combout(\Mux14~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~16 .lut_mask = 16'hADA8;
defparam \Mux14~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N14
cycloneive_lcell_comb \Mux14~17 (
// Equation(s):
// \Mux14~17_combout  = (instruction_D[21] & ((\rfile[13][17]~q ) # ((instruction_D[22])))) # (!instruction_D[21] & (((\rfile[12][17]~q  & !instruction_D[22]))))

	.dataa(\rfile[13][17]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[12][17]~q ),
	.datad(instruction_D_22),
	.cin(gnd),
	.combout(\Mux14~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~17 .lut_mask = 16'hCCB8;
defparam \Mux14~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N28
cycloneive_lcell_comb \Mux14~18 (
// Equation(s):
// \Mux14~18_combout  = (instruction_D[22] & ((\Mux14~17_combout  & ((\rfile[15][17]~q ))) # (!\Mux14~17_combout  & (\rfile[14][17]~q )))) # (!instruction_D[22] & (((\Mux14~17_combout ))))

	.dataa(\rfile[14][17]~q ),
	.datab(instruction_D_22),
	.datac(\rfile[15][17]~q ),
	.datad(\Mux14~17_combout ),
	.cin(gnd),
	.combout(\Mux14~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~18 .lut_mask = 16'hF388;
defparam \Mux14~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N2
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[25][0]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[17][0]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[17][0]~q ),
	.datad(\rfile[25][0]~q ),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hBA98;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N10
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (\Mux31~0_combout  & (((\rfile[29][0]~q )) # (!instruction_D[23]))) # (!\Mux31~0_combout  & (instruction_D[23] & ((\rfile[21][0]~q ))))

	.dataa(\Mux31~0_combout ),
	.datab(instruction_D_23),
	.datac(\rfile[29][0]~q ),
	.datad(\rfile[21][0]~q ),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hE6A2;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N6
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\rfile[27][0]~q )))) # (!instruction_D[24] & (!instruction_D[23] & (\rfile[19][0]~q )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[19][0]~q ),
	.datad(\rfile[27][0]~q ),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'hBA98;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y31_N8
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (instruction_D[23] & ((\Mux31~7_combout  & ((\rfile[31][0]~q ))) # (!\Mux31~7_combout  & (\rfile[23][0]~q )))) # (!instruction_D[23] & (\Mux31~7_combout ))

	.dataa(instruction_D_23),
	.datab(\Mux31~7_combout ),
	.datac(\rfile[23][0]~q ),
	.datad(\rfile[31][0]~q ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'hEC64;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X76_Y31_N0
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (instruction_D[23] & ((\rfile[20][0]~q ) # ((instruction_D[24])))) # (!instruction_D[23] & (((\rfile[16][0]~q  & !instruction_D[24]))))

	.dataa(\rfile[20][0]~q ),
	.datab(instruction_D_23),
	.datac(\rfile[16][0]~q ),
	.datad(instruction_D_24),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'hCCB8;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X75_Y31_N11
dffeas \rfile[28][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[28][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[28][0] .is_wysiwyg = "true";
defparam \rfile[28][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N10
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (instruction_D[24] & ((\Mux31~4_combout  & (\rfile[28][0]~q )) # (!\Mux31~4_combout  & ((\rfile[24][0]~q ))))) # (!instruction_D[24] & (\Mux31~4_combout ))

	.dataa(instruction_D_24),
	.datab(\Mux31~4_combout ),
	.datac(\rfile[28][0]~q ),
	.datad(\rfile[24][0]~q ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hE6C4;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y34_N2
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (instruction_D[24] & (instruction_D[23])) # (!instruction_D[24] & ((instruction_D[23] & (\rfile[22][0]~q )) # (!instruction_D[23] & ((\rfile[18][0]~q )))))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\rfile[22][0]~q ),
	.datad(\rfile[18][0]~q ),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hD9C8;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X74_Y34_N6
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (instruction_D[24] & ((\Mux31~2_combout  & (\rfile[30][0]~q )) # (!\Mux31~2_combout  & ((\rfile[26][0]~q ))))) # (!instruction_D[24] & (((\Mux31~2_combout ))))

	.dataa(instruction_D_24),
	.datab(\rfile[30][0]~q ),
	.datac(\rfile[26][0]~q ),
	.datad(\Mux31~2_combout ),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'hDDA0;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N28
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\Mux31~3_combout )))) # (!instruction_D[22] & (!instruction_D[21] & (\Mux31~5_combout )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\Mux31~5_combout ),
	.datad(\Mux31~3_combout ),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hBA98;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N14
cycloneive_lcell_comb \Mux31~10 (
// Equation(s):
// \Mux31~10_combout  = (instruction_D[21] & ((instruction_D[22]) # ((\rfile[5][0]~q )))) # (!instruction_D[21] & (!instruction_D[22] & (\rfile[4][0]~q )))

	.dataa(instruction_D_21),
	.datab(instruction_D_22),
	.datac(\rfile[4][0]~q ),
	.datad(\rfile[5][0]~q ),
	.cin(gnd),
	.combout(\Mux31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~10 .lut_mask = 16'hBA98;
defparam \Mux31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N30
cycloneive_lcell_comb \Mux31~11 (
// Equation(s):
// \Mux31~11_combout  = (instruction_D[22] & ((\Mux31~10_combout  & (\rfile[7][0]~q )) # (!\Mux31~10_combout  & ((\rfile[6][0]~q ))))) # (!instruction_D[22] & (\Mux31~10_combout ))

	.dataa(instruction_D_22),
	.datab(\Mux31~10_combout ),
	.datac(\rfile[7][0]~q ),
	.datad(\rfile[6][0]~q ),
	.cin(gnd),
	.combout(\Mux31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~11 .lut_mask = 16'hE6C4;
defparam \Mux31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N23
dffeas \rfile[12][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat_WB_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\rfile[12][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \rfile[12][0] .is_wysiwyg = "true";
defparam \rfile[12][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N22
cycloneive_lcell_comb \Mux31~17 (
// Equation(s):
// \Mux31~17_combout  = (instruction_D[22] & (instruction_D[21])) # (!instruction_D[22] & ((instruction_D[21] & ((\rfile[13][0]~q ))) # (!instruction_D[21] & (\rfile[12][0]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[12][0]~q ),
	.datad(\rfile[13][0]~q ),
	.cin(gnd),
	.combout(\Mux31~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~17 .lut_mask = 16'hDC98;
defparam \Mux31~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N12
cycloneive_lcell_comb \Mux31~18 (
// Equation(s):
// \Mux31~18_combout  = (instruction_D[22] & ((\Mux31~17_combout  & ((\rfile[15][0]~q ))) # (!\Mux31~17_combout  & (\rfile[14][0]~q )))) # (!instruction_D[22] & (((\Mux31~17_combout ))))

	.dataa(instruction_D_22),
	.datab(\rfile[14][0]~q ),
	.datac(\rfile[15][0]~q ),
	.datad(\Mux31~17_combout ),
	.cin(gnd),
	.combout(\Mux31~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~18 .lut_mask = 16'hF588;
defparam \Mux31~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N18
cycloneive_lcell_comb \Mux31~14 (
// Equation(s):
// \Mux31~14_combout  = (instruction_D[21] & ((instruction_D[22] & ((\rfile[3][0]~q ))) # (!instruction_D[22] & (\rfile[1][0]~q ))))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[1][0]~q ),
	.datad(\rfile[3][0]~q ),
	.cin(gnd),
	.combout(\Mux31~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~14 .lut_mask = 16'hC840;
defparam \Mux31~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N8
cycloneive_lcell_comb \Mux31~15 (
// Equation(s):
// \Mux31~15_combout  = (\Mux31~14_combout ) # ((\rfile[2][0]~q  & (!instruction_D[21] & instruction_D[22])))

	.dataa(\rfile[2][0]~q ),
	.datab(instruction_D_21),
	.datac(instruction_D_22),
	.datad(\Mux31~14_combout ),
	.cin(gnd),
	.combout(\Mux31~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~15 .lut_mask = 16'hFF20;
defparam \Mux31~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N14
cycloneive_lcell_comb \Mux31~12 (
// Equation(s):
// \Mux31~12_combout  = (instruction_D[22] & ((instruction_D[21]) # ((\rfile[10][0]~q )))) # (!instruction_D[22] & (!instruction_D[21] & (\rfile[8][0]~q )))

	.dataa(instruction_D_22),
	.datab(instruction_D_21),
	.datac(\rfile[8][0]~q ),
	.datad(\rfile[10][0]~q ),
	.cin(gnd),
	.combout(\Mux31~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~12 .lut_mask = 16'hBA98;
defparam \Mux31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N4
cycloneive_lcell_comb \Mux31~13 (
// Equation(s):
// \Mux31~13_combout  = (instruction_D[21] & ((\Mux31~12_combout  & ((\rfile[11][0]~q ))) # (!\Mux31~12_combout  & (\rfile[9][0]~q )))) # (!instruction_D[21] & (((\Mux31~12_combout ))))

	.dataa(\rfile[9][0]~q ),
	.datab(instruction_D_21),
	.datac(\rfile[11][0]~q ),
	.datad(\Mux31~12_combout ),
	.cin(gnd),
	.combout(\Mux31~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~13 .lut_mask = 16'hF388;
defparam \Mux31~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N2
cycloneive_lcell_comb \Mux31~16 (
// Equation(s):
// \Mux31~16_combout  = (instruction_D[24] & ((instruction_D[23]) # ((\Mux31~13_combout )))) # (!instruction_D[24] & (!instruction_D[23] & (\Mux31~15_combout )))

	.dataa(instruction_D_24),
	.datab(instruction_D_23),
	.datac(\Mux31~15_combout ),
	.datad(\Mux31~13_combout ),
	.cin(gnd),
	.combout(\Mux31~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~16 .lut_mask = 16'hBA98;
defparam \Mux31~16 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module memory_control (
	LessThan1,
	always0,
	dhit,
	iwait,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	LessThan1;
input 	always0;
input 	dhit;
output 	iwait;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X57_Y38_N10
cycloneive_lcell_comb \iwait~0 (
// Equation(s):
// iwait = (!dhit & (((LessThan1 & always0)) # (!\nRST~input_o )))

	.dataa(dhit),
	.datab(LessThan1),
	.datac(nRST),
	.datad(always0),
	.cin(gnd),
	.combout(iwait),
	.cout());
// synopsys translate_off
defparam \iwait~0 .lut_mask = 16'h4505;
defparam \iwait~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ram (
	is_in_use_reg,
	LessThan1,
	\ramif.ramaddr ,
	ramaddr,
	ramaddr1,
	ramaddr2,
	ramaddr3,
	ramaddr4,
	ramaddr5,
	ramaddr6,
	ramaddr7,
	ramaddr8,
	ramaddr9,
	ramaddr10,
	ramaddr11,
	ramaddr12,
	ramaddr13,
	ramaddr14,
	ramaddr15,
	ramaddr16,
	ramaddr17,
	ramWEN,
	\ramif.ramREN ,
	always0,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramstore,
	ramstore1,
	ramstore2,
	ramstore3,
	ramstore4,
	ramstore5,
	ramstore6,
	ramstore7,
	ramstore8,
	ramstore9,
	ramstore10,
	ramstore11,
	ramstore12,
	ramstore13,
	ramstore14,
	ramstore15,
	ramstore16,
	ramstore17,
	ramstore18,
	ramstore19,
	ramstore20,
	ramstore21,
	ramstore22,
	ramstore23,
	ramstore24,
	ramstore25,
	ramstore26,
	ramstore27,
	ramstore28,
	ramstore29,
	ramstore30,
	ramstore31,
	ramaddr18,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	nRST,
	nRST1,
	altera_internal_jtag1,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	is_in_use_reg;
output 	LessThan1;
input 	[31:0] \ramif.ramaddr ;
input 	ramaddr;
input 	ramaddr1;
input 	ramaddr2;
input 	ramaddr3;
input 	ramaddr4;
input 	ramaddr5;
input 	ramaddr6;
input 	ramaddr7;
input 	ramaddr8;
input 	ramaddr9;
input 	ramaddr10;
input 	ramaddr11;
input 	ramaddr12;
input 	ramaddr13;
input 	ramaddr14;
input 	ramaddr15;
input 	ramaddr16;
input 	ramaddr17;
input 	ramWEN;
input 	\ramif.ramREN ;
output 	always0;
output 	always1;
output 	ramiframload_0;
output 	ramiframload_1;
output 	ramiframload_2;
output 	ramiframload_3;
output 	ramiframload_4;
output 	ramiframload_5;
output 	ramiframload_6;
output 	ramiframload_7;
output 	ramiframload_8;
output 	ramiframload_9;
output 	ramiframload_10;
output 	ramiframload_11;
output 	ramiframload_12;
output 	ramiframload_13;
output 	ramiframload_14;
output 	ramiframload_15;
output 	ramiframload_16;
output 	ramiframload_17;
output 	ramiframload_18;
output 	ramiframload_19;
output 	ramiframload_20;
output 	ramiframload_21;
output 	ramiframload_22;
output 	ramiframload_23;
output 	ramiframload_24;
output 	ramiframload_25;
output 	ramiframload_26;
output 	ramiframload_27;
output 	ramiframload_28;
output 	ramiframload_29;
output 	ramiframload_30;
output 	ramiframload_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramstore;
input 	ramstore1;
input 	ramstore2;
input 	ramstore3;
input 	ramstore4;
input 	ramstore5;
input 	ramstore6;
input 	ramstore7;
input 	ramstore8;
input 	ramstore9;
input 	ramstore10;
input 	ramstore11;
input 	ramstore12;
input 	ramstore13;
input 	ramstore14;
input 	ramstore15;
input 	ramstore16;
input 	ramstore17;
input 	ramstore18;
input 	ramstore19;
input 	ramstore20;
input 	ramstore21;
input 	ramstore22;
input 	ramstore23;
input 	ramstore24;
input 	ramstore25;
input 	ramstore26;
input 	ramstore27;
input 	ramstore28;
input 	ramstore29;
input 	ramstore30;
input 	ramstore31;
input 	ramaddr18;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	nRST;
input 	nRST1;
input 	altera_internal_jtag1;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ;
wire \always0~2_combout ;
wire \always0~5_combout ;
wire \always0~12_combout ;
wire \always0~15_combout ;
wire \Add0~0_combout ;
wire \addr[22]~feeder_combout ;
wire \addr[25]~feeder_combout ;
wire \addr[24]~feeder_combout ;
wire \always0~0_combout ;
wire \addr[2]~feeder_combout ;
wire \always0~1_combout ;
wire \addr[6]~feeder_combout ;
wire \always0~3_combout ;
wire \always0~4_combout ;
wire \always0~22_combout ;
wire \always0~8_combout ;
wire \always0~6_combout ;
wire \always0~7_combout ;
wire \always0~9_combout ;
wire \always0~23_combout ;
wire \count[2]~1_combout ;
wire \count[0]~3_combout ;
wire \count[3]~0_combout ;
wire \count[1]~2_combout ;
wire \always0~16_combout ;
wire \always0~18_combout ;
wire \always0~17_combout ;
wire \always0~19_combout ;
wire \always0~11_combout ;
wire \always0~13_combout ;
wire \always0~10_combout ;
wire \always0~14_combout ;
wire \always0~20_combout ;
wire [1:0] en;
wire [3:0] count;
wire [31:0] addr;
wire [0:0] \altsyncram_component|auto_generated|altsyncram1|address_reg_a ;


altsyncram_1 altsyncram_component(
	.ram_block3a32(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.ram_block3a0(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.ram_block3a33(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.ram_block3a1(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.ram_block3a34(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.ram_block3a2(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.ram_block3a35(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.ram_block3a3(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.ram_block3a36(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.ram_block3a4(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.ram_block3a37(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.ram_block3a5(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.ram_block3a38(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.ram_block3a6(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.ram_block3a39(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.ram_block3a7(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.ram_block3a40(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.ram_block3a8(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.ram_block3a41(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.ram_block3a9(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.ram_block3a42(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.ram_block3a10(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.ram_block3a43(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.ram_block3a11(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.ram_block3a44(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.ram_block3a12(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.ram_block3a45(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.ram_block3a13(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.ram_block3a46(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.ram_block3a14(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.ram_block3a47(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.ram_block3a15(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.ram_block3a48(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.ram_block3a16(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.ram_block3a49(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.ram_block3a17(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.ram_block3a50(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.ram_block3a18(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.ram_block3a51(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.ram_block3a19(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.ram_block3a52(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.ram_block3a20(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.ram_block3a53(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.ram_block3a21(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.ram_block3a54(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.ram_block3a22(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.ram_block3a55(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.ram_block3a23(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.ram_block3a56(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.ram_block3a24(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.ram_block3a57(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.ram_block3a25(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.ram_block3a58(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.ram_block3a26(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.ram_block3a59(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.ram_block3a27(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.ram_block3a60(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.ram_block3a28(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.ram_block3a61(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.ram_block3a29(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.ram_block3a62(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.ram_block3a30(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.ram_block3a63(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.ram_block3a31(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.address_a({gnd,ramaddr13,ramaddr10,ramaddr11,ramaddr8,ramaddr9,ramaddr6,ramaddr7,ramaddr4,ramaddr5,ramaddr2,ramaddr3,ramaddr,ramaddr1}),
	.ramaddr(ramaddr12),
	.ramWEN(ramWEN),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({ramstore31,ramstore30,ramstore29,ramstore28,ramstore27,ramstore26,ramstore25,ramstore24,ramstore23,ramstore22,ramstore21,ramstore20,ramstore19,ramstore18,ramstore17,ramstore16,ramstore15,ramstore14,ramstore13,ramstore12,ramstore11,ramstore10,ramstore9,ramstore8,ramstore7,ramstore6,
ramstore5,ramstore4,ramstore3,ramstore2,ramstore1,ramstore}),
	.ramaddr1(ramaddr18),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X53_Y35_N31
dffeas \addr[1] (
	.clk(CLK),
	.d(\ramif.ramaddr [1]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[1] .is_wysiwyg = "true";
defparam \addr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N17
dffeas \addr[4] (
	.clk(CLK),
	.d(ramaddr3),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[4] .is_wysiwyg = "true";
defparam \addr[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N23
dffeas \addr[5] (
	.clk(CLK),
	.d(ramaddr2),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[5] .is_wysiwyg = "true";
defparam \addr[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N10
cycloneive_lcell_comb \always0~2 (
// Equation(s):
// \always0~2_combout  = (addr[5] & (\ramaddr~9_combout  & (addr[4] $ (!\ramaddr~11_combout )))) # (!addr[5] & (!\ramaddr~9_combout  & (addr[4] $ (!\ramaddr~11_combout ))))

	.dataa(addr[5]),
	.datab(addr[4]),
	.datac(ramaddr3),
	.datad(ramaddr2),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
// synopsys translate_off
defparam \always0~2 .lut_mask = 16'h8241;
defparam \always0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N3
dffeas \addr[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr4),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[7] .is_wysiwyg = "true";
defparam \addr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N21
dffeas \addr[8] (
	.clk(CLK),
	.d(ramaddr7),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[8] .is_wysiwyg = "true";
defparam \addr[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N27
dffeas \addr[9] (
	.clk(CLK),
	.d(ramaddr6),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[9] .is_wysiwyg = "true";
defparam \addr[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N0
cycloneive_lcell_comb \always0~5 (
// Equation(s):
// \always0~5_combout  = (\ramaddr~17_combout  & (addr[9] & (addr[8] $ (!\ramaddr~19_combout )))) # (!\ramaddr~17_combout  & (!addr[9] & (addr[8] $ (!\ramaddr~19_combout ))))

	.dataa(ramaddr6),
	.datab(addr[8]),
	.datac(addr[9]),
	.datad(ramaddr7),
	.cin(gnd),
	.combout(\always0~5_combout ),
	.cout());
// synopsys translate_off
defparam \always0~5 .lut_mask = 16'h8421;
defparam \always0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N19
dffeas \addr[11] (
	.clk(CLK),
	.d(ramaddr8),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[11] .is_wysiwyg = "true";
defparam \addr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y38_N17
dffeas \addr[13] (
	.clk(CLK),
	.d(ramaddr10),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[13] .is_wysiwyg = "true";
defparam \addr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N23
dffeas \addr[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr13),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[14] .is_wysiwyg = "true";
defparam \addr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N11
dffeas \addr[16] (
	.clk(CLK),
	.d(\ramif.ramaddr [16]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[16] .is_wysiwyg = "true";
defparam \addr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N5
dffeas \addr[18] (
	.clk(CLK),
	.d(\ramif.ramaddr [18]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[18] .is_wysiwyg = "true";
defparam \addr[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N3
dffeas \addr[20] (
	.clk(CLK),
	.d(\ramif.ramaddr [20]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[20] .is_wysiwyg = "true";
defparam \addr[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N5
dffeas \addr[21] (
	.clk(CLK),
	.d(\ramif.ramaddr [21]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[21] .is_wysiwyg = "true";
defparam \addr[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N8
cycloneive_lcell_comb \always0~12 (
// Equation(s):
// \always0~12_combout  = (addr[20] & (\ramaddr~43_combout  & (\ramaddr~41_combout  $ (!addr[21])))) # (!addr[20] & (!\ramaddr~43_combout  & (\ramaddr~41_combout  $ (!addr[21]))))

	.dataa(addr[20]),
	.datab(\ramif.ramaddr [21]),
	.datac(addr[21]),
	.datad(\ramif.ramaddr [20]),
	.cin(gnd),
	.combout(\always0~12_combout ),
	.cout());
// synopsys translate_off
defparam \always0~12 .lut_mask = 16'h8241;
defparam \always0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N13
dffeas \addr[22] (
	.clk(CLK),
	.d(\addr[22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[22] .is_wysiwyg = "true";
defparam \addr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N1
dffeas \addr[24] (
	.clk(CLK),
	.d(\addr[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[24] .is_wysiwyg = "true";
defparam \addr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N7
dffeas \addr[25] (
	.clk(CLK),
	.d(\addr[25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[25] .is_wysiwyg = "true";
defparam \addr[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N18
cycloneive_lcell_comb \always0~15 (
// Equation(s):
// \always0~15_combout  = (addr[25] & (\ramaddr~49_combout  & (addr[24] $ (!\ramaddr~51_combout )))) # (!addr[25] & (!\ramaddr~49_combout  & (addr[24] $ (!\ramaddr~51_combout ))))

	.dataa(addr[25]),
	.datab(addr[24]),
	.datac(ramaddr17),
	.datad(ramaddr16),
	.cin(gnd),
	.combout(\always0~15_combout ),
	.cout());
// synopsys translate_off
defparam \always0~15 .lut_mask = 16'h8241;
defparam \always0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y36_N31
dffeas \addr[26] (
	.clk(CLK),
	.d(\ramif.ramaddr [26]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[26]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[26] .is_wysiwyg = "true";
defparam \addr[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N15
dffeas \addr[28] (
	.clk(CLK),
	.d(\ramif.ramaddr [28]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[28]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[28] .is_wysiwyg = "true";
defparam \addr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N9
dffeas \addr[31] (
	.clk(CLK),
	.d(\ramif.ramaddr [31]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[31]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[31] .is_wysiwyg = "true";
defparam \addr[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N30
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = (count[0] & count[1])

	.dataa(gnd),
	.datab(count[0]),
	.datac(gnd),
	.datad(count[1]),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'hCC00;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N12
cycloneive_lcell_comb \addr[22]~feeder (
// Equation(s):
// \addr[22]~feeder_combout  = \ramaddr~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr15),
	.cin(gnd),
	.combout(\addr[22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[22]~feeder .lut_mask = 16'hFF00;
defparam \addr[22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N6
cycloneive_lcell_comb \addr[25]~feeder (
// Equation(s):
// \addr[25]~feeder_combout  = \ramaddr~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr16),
	.cin(gnd),
	.combout(\addr[25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[25]~feeder .lut_mask = 16'hFF00;
defparam \addr[25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N0
cycloneive_lcell_comb \addr[24]~feeder (
// Equation(s):
// \addr[24]~feeder_combout  = \ramaddr~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(ramaddr17),
	.datad(gnd),
	.cin(gnd),
	.combout(\addr[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[24]~feeder .lut_mask = 16'hF0F0;
defparam \addr[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N26
cycloneive_lcell_comb \LessThan1~0 (
// Equation(s):
// LessThan1 = (count[3]) # ((count[2] & (count[0] & count[1])))

	.dataa(count[2]),
	.datab(count[0]),
	.datac(count[3]),
	.datad(count[1]),
	.cin(gnd),
	.combout(LessThan1),
	.cout());
// synopsys translate_off
defparam \LessThan1~0 .lut_mask = 16'hF8F0;
defparam \LessThan1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N24
cycloneive_lcell_comb \always0~21 (
// Equation(s):
// always0 = (\always0~9_combout  & (\always0~20_combout  & \always0~4_combout ))

	.dataa(gnd),
	.datab(\always0~9_combout ),
	.datac(\always0~20_combout ),
	.datad(\always0~4_combout ),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~21 .lut_mask = 16'hC000;
defparam \always0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N6
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// always1 = ((LessThan1 & always0)) # (!\nRST~input_o )

	.dataa(gnd),
	.datab(LessThan1),
	.datac(nRST),
	.datad(always0),
	.cin(gnd),
	.combout(always1),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'hCF0F;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N16
cycloneive_lcell_comb \ramif.ramload[0]~0 (
// Equation(s):
// ramiframload_0 = ((address_reg_a_0 & ((ram_block3a321))) # (!address_reg_a_0 & (ram_block3a01))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.cin(gnd),
	.combout(ramiframload_0),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~0 .lut_mask = 16'hFB73;
defparam \ramif.ramload[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N14
cycloneive_lcell_comb \ramif.ramload[1]~1 (
// Equation(s):
// ramiframload_1 = (always1 & ((address_reg_a_0 & ((ram_block3a331))) # (!address_reg_a_0 & (ram_block3a110))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.cin(gnd),
	.combout(ramiframload_1),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~1 .lut_mask = 16'hC808;
defparam \ramif.ramload[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N4
cycloneive_lcell_comb \ramif.ramload[2]~2 (
// Equation(s):
// ramiframload_2 = (always1 & ((address_reg_a_0 & (ram_block3a341)) # (!address_reg_a_0 & ((ram_block3a210)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_2),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[2]~2 .lut_mask = 16'hB800;
defparam \ramif.ramload[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N26
cycloneive_lcell_comb \ramif.ramload[3]~3 (
// Equation(s):
// ramiframload_3 = (always1 & ((address_reg_a_0 & (ram_block3a351)) # (!address_reg_a_0 & ((ram_block3a310)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_3),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[3]~3 .lut_mask = 16'hB800;
defparam \ramif.ramload[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N0
cycloneive_lcell_comb \ramif.ramload[4]~4 (
// Equation(s):
// ramiframload_4 = ((address_reg_a_0 & (ram_block3a361)) # (!address_reg_a_0 & ((ram_block3a410)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_4),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[4]~4 .lut_mask = 16'hACFF;
defparam \ramif.ramload[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N8
cycloneive_lcell_comb \ramif.ramload[5]~5 (
// Equation(s):
// ramiframload_5 = (always1 & ((address_reg_a_0 & ((ram_block3a371))) # (!address_reg_a_0 & (ram_block3a510))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.cin(gnd),
	.combout(ramiframload_5),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[5]~5 .lut_mask = 16'hE020;
defparam \ramif.ramload[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N26
cycloneive_lcell_comb \ramif.ramload[6]~6 (
// Equation(s):
// ramiframload_6 = ((address_reg_a_0 & (ram_block3a381)) # (!address_reg_a_0 & ((ram_block3a64)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_6),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[6]~6 .lut_mask = 16'hACFF;
defparam \ramif.ramload[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N16
cycloneive_lcell_comb \ramif.ramload[7]~7 (
// Equation(s):
// ramiframload_7 = ((address_reg_a_0 & ((ram_block3a391))) # (!address_reg_a_0 & (ram_block3a71))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_7),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[7]~7 .lut_mask = 16'hE2FF;
defparam \ramif.ramload[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N12
cycloneive_lcell_comb \ramif.ramload[8]~8 (
// Equation(s):
// ramiframload_8 = (always1 & ((address_reg_a_0 & ((ram_block3a401))) # (!address_reg_a_0 & (ram_block3a81))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_8),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[8]~8 .lut_mask = 16'hCA00;
defparam \ramif.ramload[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N16
cycloneive_lcell_comb \ramif.ramload[9]~9 (
// Equation(s):
// ramiframload_9 = ((address_reg_a_0 & ((ram_block3a412))) # (!address_reg_a_0 & (ram_block3a91))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_9),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[9]~9 .lut_mask = 16'hE2FF;
defparam \ramif.ramload[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N10
cycloneive_lcell_comb \ramif.ramload[10]~10 (
// Equation(s):
// ramiframload_10 = (always1 & ((address_reg_a_0 & ((ram_block3a421))) # (!address_reg_a_0 & (ram_block3a101))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_10),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[10]~10 .lut_mask = 16'hCA00;
defparam \ramif.ramload[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N24
cycloneive_lcell_comb \ramif.ramload[11]~11 (
// Equation(s):
// ramiframload_11 = ((address_reg_a_0 & ((ram_block3a431))) # (!address_reg_a_0 & (ram_block3a112))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_11),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[11]~11 .lut_mask = 16'hE2FF;
defparam \ramif.ramload[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N16
cycloneive_lcell_comb \ramif.ramload[12]~12 (
// Equation(s):
// ramiframload_12 = ((address_reg_a_0 & (ram_block3a441)) # (!address_reg_a_0 & ((ram_block3a121)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_12),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[12]~12 .lut_mask = 16'hDDF5;
defparam \ramif.ramload[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N2
cycloneive_lcell_comb \ramif.ramload[13]~13 (
// Equation(s):
// ramiframload_13 = ((address_reg_a_0 & ((ram_block3a451))) # (!address_reg_a_0 & (ram_block3a131))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_13),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[13]~13 .lut_mask = 16'hE2FF;
defparam \ramif.ramload[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N22
cycloneive_lcell_comb \ramif.ramload[14]~14 (
// Equation(s):
// ramiframload_14 = (always1 & ((address_reg_a_0 & ((ram_block3a461))) # (!address_reg_a_0 & (ram_block3a141))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_14),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[14]~14 .lut_mask = 16'hE200;
defparam \ramif.ramload[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N24
cycloneive_lcell_comb \ramif.ramload[15]~15 (
// Equation(s):
// ramiframload_15 = ((address_reg_a_0 & ((ram_block3a471))) # (!address_reg_a_0 & (ram_block3a151))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.cin(gnd),
	.combout(ramiframload_15),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[15]~15 .lut_mask = 16'hFD5D;
defparam \ramif.ramload[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N16
cycloneive_lcell_comb \ramif.ramload[16]~16 (
// Equation(s):
// ramiframload_16 = ((address_reg_a_0 & ((ram_block3a481))) # (!address_reg_a_0 & (ram_block3a161))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_16),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~16 .lut_mask = 16'hE4FF;
defparam \ramif.ramload[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N8
cycloneive_lcell_comb \ramif.ramload[17]~17 (
// Equation(s):
// ramiframload_17 = (always1 & ((address_reg_a_0 & (ram_block3a491)) # (!address_reg_a_0 & ((ram_block3a171)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_17),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~17 .lut_mask = 16'hD800;
defparam \ramif.ramload[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N20
cycloneive_lcell_comb \ramif.ramload[18]~18 (
// Equation(s):
// ramiframload_18 = (always1 & ((address_reg_a_0 & (ram_block3a501)) # (!address_reg_a_0 & ((ram_block3a181)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_18),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[18]~18 .lut_mask = 16'hB800;
defparam \ramif.ramload[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N18
cycloneive_lcell_comb \ramif.ramload[19]~19 (
// Equation(s):
// ramiframload_19 = (always1 & ((address_reg_a_0 & (ram_block3a512)) # (!address_reg_a_0 & ((ram_block3a191)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_19),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[19]~19 .lut_mask = 16'hB800;
defparam \ramif.ramload[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N8
cycloneive_lcell_comb \ramif.ramload[20]~20 (
// Equation(s):
// ramiframload_20 = ((address_reg_a_0 & ((ram_block3a521))) # (!address_reg_a_0 & (ram_block3a201))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_20),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[20]~20 .lut_mask = 16'hCAFF;
defparam \ramif.ramload[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N10
cycloneive_lcell_comb \ramif.ramload[21]~21 (
// Equation(s):
// ramiframload_21 = (always1 & ((address_reg_a_0 & ((ram_block3a531))) # (!address_reg_a_0 & (ram_block3a212))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.cin(gnd),
	.combout(ramiframload_21),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[21]~21 .lut_mask = 16'hC840;
defparam \ramif.ramload[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N16
cycloneive_lcell_comb \ramif.ramload[22]~22 (
// Equation(s):
// ramiframload_22 = ((address_reg_a_0 & (ram_block3a541)) # (!address_reg_a_0 & ((ram_block3a221)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.cin(gnd),
	.combout(ramiframload_22),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[22]~22 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N24
cycloneive_lcell_comb \ramif.ramload[23]~23 (
// Equation(s):
// ramiframload_23 = ((address_reg_a_0 & ((ram_block3a551))) # (!address_reg_a_0 & (ram_block3a231))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_23),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[23]~23 .lut_mask = 16'hE2FF;
defparam \ramif.ramload[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N14
cycloneive_lcell_comb \ramif.ramload[24]~24 (
// Equation(s):
// ramiframload_24 = (always1 & ((address_reg_a_0 & (ram_block3a561)) # (!address_reg_a_0 & ((ram_block3a241)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_24),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[24]~24 .lut_mask = 16'hAC00;
defparam \ramif.ramload[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N8
cycloneive_lcell_comb \ramif.ramload[25]~25 (
// Equation(s):
// ramiframload_25 = ((address_reg_a_0 & (ram_block3a571)) # (!address_reg_a_0 & ((ram_block3a251)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_25),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[25]~25 .lut_mask = 16'hB8FF;
defparam \ramif.ramload[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N28
cycloneive_lcell_comb \ramif.ramload[26]~26 (
// Equation(s):
// ramiframload_26 = (always1 & ((address_reg_a_0 & ((ram_block3a581))) # (!address_reg_a_0 & (ram_block3a261))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.cin(gnd),
	.combout(ramiframload_26),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~26 .lut_mask = 16'hA820;
defparam \ramif.ramload[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N20
cycloneive_lcell_comb \ramif.ramload[27]~27 (
// Equation(s):
// ramiframload_27 = ((address_reg_a_0 & ((ram_block3a591))) # (!address_reg_a_0 & (ram_block3a271))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.cin(gnd),
	.combout(ramiframload_27),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~27 .lut_mask = 16'hEF4F;
defparam \ramif.ramload[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N22
cycloneive_lcell_comb \ramif.ramload[28]~28 (
// Equation(s):
// ramiframload_28 = ((address_reg_a_0 & ((ram_block3a601))) # (!address_reg_a_0 & (ram_block3a281))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.cin(gnd),
	.combout(ramiframload_28),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~28 .lut_mask = 16'hEF4F;
defparam \ramif.ramload[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N0
cycloneive_lcell_comb \ramif.ramload[29]~29 (
// Equation(s):
// ramiframload_29 = ((address_reg_a_0 & (ram_block3a611)) # (!address_reg_a_0 & ((ram_block3a291)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_29),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~29 .lut_mask = 16'hACFF;
defparam \ramif.ramload[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N10
cycloneive_lcell_comb \ramif.ramload[30]~30 (
// Equation(s):
// ramiframload_30 = (always1 & ((address_reg_a_0 & (ram_block3a621)) # (!address_reg_a_0 & ((ram_block3a301)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_30),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~30 .lut_mask = 16'hD800;
defparam \ramif.ramload[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N8
cycloneive_lcell_comb \ramif.ramload[31]~31 (
// Equation(s):
// ramiframload_31 = ((address_reg_a_0 & ((ram_block3a631))) # (!address_reg_a_0 & (ram_block3a312))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_31),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~31 .lut_mask = 16'hCAFF;
defparam \ramif.ramload[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N21
dffeas \addr[0] (
	.clk(CLK),
	.d(\ramif.ramaddr [0]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[0] .is_wysiwyg = "true";
defparam \addr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N14
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (addr[1] & (\ramaddr~1_combout  & (addr[0] $ (!\ramaddr~3_combout )))) # (!addr[1] & (!\ramaddr~1_combout  & (addr[0] $ (!\ramaddr~3_combout ))))

	.dataa(addr[1]),
	.datab(addr[0]),
	.datac(\ramif.ramaddr [0]),
	.datad(\ramif.ramaddr [1]),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h8241;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N1
dffeas \addr[3] (
	.clk(CLK),
	.d(ramaddr),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[3] .is_wysiwyg = "true";
defparam \addr[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N12
cycloneive_lcell_comb \addr[2]~feeder (
// Equation(s):
// \addr[2]~feeder_combout  = \ramaddr~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr1),
	.cin(gnd),
	.combout(\addr[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[2]~feeder .lut_mask = 16'hFF00;
defparam \addr[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N13
dffeas \addr[2] (
	.clk(CLK),
	.d(\addr[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[2] .is_wysiwyg = "true";
defparam \addr[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N20
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = (\ramaddr~5_combout  & (addr[3] & (addr[2] $ (!\ramaddr~7_combout )))) # (!\ramaddr~5_combout  & (!addr[3] & (addr[2] $ (!\ramaddr~7_combout ))))

	.dataa(ramaddr),
	.datab(addr[3]),
	.datac(addr[2]),
	.datad(ramaddr1),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'h9009;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N22
cycloneive_lcell_comb \addr[6]~feeder (
// Equation(s):
// \addr[6]~feeder_combout  = \ramaddr~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr5),
	.cin(gnd),
	.combout(\addr[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[6]~feeder .lut_mask = 16'hFF00;
defparam \addr[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y36_N23
dffeas \addr[6] (
	.clk(CLK),
	.d(\addr[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[6] .is_wysiwyg = "true";
defparam \addr[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N18
cycloneive_lcell_comb \always0~3 (
// Equation(s):
// \always0~3_combout  = (addr[7] & (\ramaddr~13_combout  & (\ramaddr~15_combout  $ (!addr[6])))) # (!addr[7] & (!\ramaddr~13_combout  & (\ramaddr~15_combout  $ (!addr[6]))))

	.dataa(addr[7]),
	.datab(ramaddr5),
	.datac(addr[6]),
	.datad(ramaddr4),
	.cin(gnd),
	.combout(\always0~3_combout ),
	.cout());
// synopsys translate_off
defparam \always0~3 .lut_mask = 16'h8241;
defparam \always0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N0
cycloneive_lcell_comb \always0~4 (
// Equation(s):
// \always0~4_combout  = (\always0~2_combout  & (\always0~0_combout  & (\always0~1_combout  & \always0~3_combout )))

	.dataa(\always0~2_combout ),
	.datab(\always0~0_combout ),
	.datac(\always0~1_combout ),
	.datad(\always0~3_combout ),
	.cin(gnd),
	.combout(\always0~4_combout ),
	.cout());
// synopsys translate_off
defparam \always0~4 .lut_mask = 16'h8000;
defparam \always0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N27
dffeas \en[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramWEN),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[0]),
	.prn(vcc));
// synopsys translate_off
defparam \en[0] .is_wysiwyg = "true";
defparam \en[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N13
dffeas \en[1] (
	.clk(CLK),
	.d(\ramif.ramREN ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[1]),
	.prn(vcc));
// synopsys translate_off
defparam \en[1] .is_wysiwyg = "true";
defparam \en[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N26
cycloneive_lcell_comb \always0~22 (
// Equation(s):
// \always0~22_combout  = (\ramREN~0_combout  & ((\ramWEN~0_combout  $ (en[0])) # (!en[1]))) # (!\ramREN~0_combout  & ((en[1]) # (\ramWEN~0_combout  $ (en[0]))))

	.dataa(\ramif.ramREN ),
	.datab(ramWEN),
	.datac(en[0]),
	.datad(en[1]),
	.cin(gnd),
	.combout(\always0~22_combout ),
	.cout());
// synopsys translate_off
defparam \always0~22 .lut_mask = 16'h7DBE;
defparam \always0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y38_N5
dffeas \addr[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr18),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[15] .is_wysiwyg = "true";
defparam \addr[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N4
cycloneive_lcell_comb \always0~8 (
// Equation(s):
// \always0~8_combout  = (addr[14] & (\ramaddr~31_combout  & (addr[15] $ (\ramaddr~29_combout )))) # (!addr[14] & (!\ramaddr~31_combout  & (addr[15] $ (\ramaddr~29_combout ))))

	.dataa(addr[14]),
	.datab(ramaddr13),
	.datac(addr[15]),
	.datad(ramaddr12),
	.cin(gnd),
	.combout(\always0~8_combout ),
	.cout());
// synopsys translate_off
defparam \always0~8 .lut_mask = 16'h0990;
defparam \always0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N25
dffeas \addr[10] (
	.clk(CLK),
	.d(ramaddr9),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[10] .is_wysiwyg = "true";
defparam \addr[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N8
cycloneive_lcell_comb \always0~6 (
// Equation(s):
// \always0~6_combout  = (addr[11] & (\ramaddr~21_combout  & (addr[10] $ (!\ramaddr~23_combout )))) # (!addr[11] & (!\ramaddr~21_combout  & (addr[10] $ (!\ramaddr~23_combout ))))

	.dataa(addr[11]),
	.datab(addr[10]),
	.datac(ramaddr9),
	.datad(ramaddr8),
	.cin(gnd),
	.combout(\always0~6_combout ),
	.cout());
// synopsys translate_off
defparam \always0~6 .lut_mask = 16'h8241;
defparam \always0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N7
dffeas \addr[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr11),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[12] .is_wysiwyg = "true";
defparam \addr[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N6
cycloneive_lcell_comb \always0~7 (
// Equation(s):
// \always0~7_combout  = (addr[13] & (\ramaddr~25_combout  & (addr[12] $ (!\ramaddr~27_combout )))) # (!addr[13] & (!\ramaddr~25_combout  & (addr[12] $ (!\ramaddr~27_combout ))))

	.dataa(addr[13]),
	.datab(ramaddr10),
	.datac(addr[12]),
	.datad(ramaddr11),
	.cin(gnd),
	.combout(\always0~7_combout ),
	.cout());
// synopsys translate_off
defparam \always0~7 .lut_mask = 16'h9009;
defparam \always0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N2
cycloneive_lcell_comb \always0~9 (
// Equation(s):
// \always0~9_combout  = (\always0~5_combout  & (\always0~8_combout  & (\always0~6_combout  & \always0~7_combout )))

	.dataa(\always0~5_combout ),
	.datab(\always0~8_combout ),
	.datac(\always0~6_combout ),
	.datad(\always0~7_combout ),
	.cin(gnd),
	.combout(\always0~9_combout ),
	.cout());
// synopsys translate_off
defparam \always0~9 .lut_mask = 16'h8000;
defparam \always0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N20
cycloneive_lcell_comb \always0~23 (
// Equation(s):
// \always0~23_combout  = (((\always0~22_combout ) # (!\always0~9_combout )) # (!\always0~4_combout )) # (!\always0~20_combout )

	.dataa(\always0~20_combout ),
	.datab(\always0~4_combout ),
	.datac(\always0~22_combout ),
	.datad(\always0~9_combout ),
	.cin(gnd),
	.combout(\always0~23_combout ),
	.cout());
// synopsys translate_off
defparam \always0~23 .lut_mask = 16'hF7FF;
defparam \always0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N10
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = (!\always0~23_combout  & (count[2] $ (((\Add0~0_combout  & !LessThan1)))))

	.dataa(\Add0~0_combout ),
	.datab(\always0~23_combout ),
	.datac(count[2]),
	.datad(LessThan1),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h3012;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N11
dffeas \count[2] (
	.clk(CLK),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N30
cycloneive_lcell_comb \count[0]~3 (
// Equation(s):
// \count[0]~3_combout  = (!\always0~23_combout  & (LessThan1 $ (!count[0])))

	.dataa(gnd),
	.datab(LessThan1),
	.datac(count[0]),
	.datad(\always0~23_combout ),
	.cin(gnd),
	.combout(\count[0]~3_combout ),
	.cout());
// synopsys translate_off
defparam \count[0]~3 .lut_mask = 16'h00C3;
defparam \count[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N31
dffeas \count[0] (
	.clk(CLK),
	.d(\count[0]~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N4
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = (!\always0~23_combout  & count[3])

	.dataa(gnd),
	.datab(\always0~23_combout ),
	.datac(count[3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h3030;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N5
dffeas \count[3] (
	.clk(CLK),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N12
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = (!\always0~23_combout  & (count[1] $ (((count[0] & !LessThan1)))))

	.dataa(count[0]),
	.datab(LessThan1),
	.datac(count[1]),
	.datad(\always0~23_combout ),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h00D2;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N13
dffeas \count[1] (
	.clk(CLK),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N9
dffeas \addr[27] (
	.clk(CLK),
	.d(\ramif.ramaddr [27]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[27]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[27] .is_wysiwyg = "true";
defparam \addr[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N14
cycloneive_lcell_comb \always0~16 (
// Equation(s):
// \always0~16_combout  = (addr[26] & (\ramaddr~55_combout  & (addr[27] $ (!\ramaddr~53_combout )))) # (!addr[26] & (!\ramaddr~55_combout  & (addr[27] $ (!\ramaddr~53_combout ))))

	.dataa(addr[26]),
	.datab(addr[27]),
	.datac(\ramif.ramaddr [26]),
	.datad(\ramif.ramaddr [27]),
	.cin(gnd),
	.combout(\always0~16_combout ),
	.cout());
// synopsys translate_off
defparam \always0~16 .lut_mask = 16'h8421;
defparam \always0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N19
dffeas \addr[30] (
	.clk(CLK),
	.d(\ramif.ramaddr [30]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[30]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[30] .is_wysiwyg = "true";
defparam \addr[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N14
cycloneive_lcell_comb \always0~18 (
// Equation(s):
// \always0~18_combout  = (addr[31] & (\ramaddr~61_combout  & (addr[30] $ (!\ramaddr~63_combout )))) # (!addr[31] & (!\ramaddr~61_combout  & (addr[30] $ (!\ramaddr~63_combout ))))

	.dataa(addr[31]),
	.datab(addr[30]),
	.datac(\ramif.ramaddr [31]),
	.datad(\ramif.ramaddr [30]),
	.cin(gnd),
	.combout(\always0~18_combout ),
	.cout());
// synopsys translate_off
defparam \always0~18 .lut_mask = 16'h8421;
defparam \always0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N25
dffeas \addr[29] (
	.clk(CLK),
	.d(\ramif.ramaddr [29]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[29]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[29] .is_wysiwyg = "true";
defparam \addr[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N30
cycloneive_lcell_comb \always0~17 (
// Equation(s):
// \always0~17_combout  = (addr[28] & (\ramaddr~59_combout  & (addr[29] $ (!\ramaddr~57_combout )))) # (!addr[28] & (!\ramaddr~59_combout  & (addr[29] $ (!\ramaddr~57_combout ))))

	.dataa(addr[28]),
	.datab(addr[29]),
	.datac(\ramif.ramaddr [28]),
	.datad(\ramif.ramaddr [29]),
	.cin(gnd),
	.combout(\always0~17_combout ),
	.cout());
// synopsys translate_off
defparam \always0~17 .lut_mask = 16'h8421;
defparam \always0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N14
cycloneive_lcell_comb \always0~19 (
// Equation(s):
// \always0~19_combout  = (\always0~15_combout  & (\always0~16_combout  & (\always0~18_combout  & \always0~17_combout )))

	.dataa(\always0~15_combout ),
	.datab(\always0~16_combout ),
	.datac(\always0~18_combout ),
	.datad(\always0~17_combout ),
	.cin(gnd),
	.combout(\always0~19_combout ),
	.cout());
// synopsys translate_off
defparam \always0~19 .lut_mask = 16'h8000;
defparam \always0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N3
dffeas \addr[19] (
	.clk(CLK),
	.d(\ramif.ramaddr [19]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[19] .is_wysiwyg = "true";
defparam \addr[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N26
cycloneive_lcell_comb \always0~11 (
// Equation(s):
// \always0~11_combout  = (addr[18] & (\ramaddr~39_combout  & (addr[19] $ (!\ramaddr~37_combout )))) # (!addr[18] & (!\ramaddr~39_combout  & (addr[19] $ (!\ramaddr~37_combout ))))

	.dataa(addr[18]),
	.datab(addr[19]),
	.datac(\ramif.ramaddr [18]),
	.datad(\ramif.ramaddr [19]),
	.cin(gnd),
	.combout(\always0~11_combout ),
	.cout());
// synopsys translate_off
defparam \always0~11 .lut_mask = 16'h8421;
defparam \always0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N27
dffeas \addr[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr14),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[23] .is_wysiwyg = "true";
defparam \addr[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N26
cycloneive_lcell_comb \always0~13 (
// Equation(s):
// \always0~13_combout  = (addr[22] & (\ramaddr~47_combout  & (\ramaddr~45_combout  $ (!addr[23])))) # (!addr[22] & (!\ramaddr~47_combout  & (\ramaddr~45_combout  $ (!addr[23]))))

	.dataa(addr[22]),
	.datab(ramaddr14),
	.datac(addr[23]),
	.datad(ramaddr15),
	.cin(gnd),
	.combout(\always0~13_combout ),
	.cout());
// synopsys translate_off
defparam \always0~13 .lut_mask = 16'h8241;
defparam \always0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y36_N25
dffeas \addr[17] (
	.clk(CLK),
	.d(\ramif.ramaddr [17]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[17] .is_wysiwyg = "true";
defparam \addr[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N12
cycloneive_lcell_comb \always0~10 (
// Equation(s):
// \always0~10_combout  = (addr[16] & (\ramaddr~35_combout  & (addr[17] $ (!\ramaddr~33_combout )))) # (!addr[16] & (!\ramaddr~35_combout  & (addr[17] $ (!\ramaddr~33_combout ))))

	.dataa(addr[16]),
	.datab(addr[17]),
	.datac(\ramif.ramaddr [16]),
	.datad(\ramif.ramaddr [17]),
	.cin(gnd),
	.combout(\always0~10_combout ),
	.cout());
// synopsys translate_off
defparam \always0~10 .lut_mask = 16'h8421;
defparam \always0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N16
cycloneive_lcell_comb \always0~14 (
// Equation(s):
// \always0~14_combout  = (\always0~12_combout  & (\always0~11_combout  & (\always0~13_combout  & \always0~10_combout )))

	.dataa(\always0~12_combout ),
	.datab(\always0~11_combout ),
	.datac(\always0~13_combout ),
	.datad(\always0~10_combout ),
	.cin(gnd),
	.combout(\always0~14_combout ),
	.cout());
// synopsys translate_off
defparam \always0~14 .lut_mask = 16'h8000;
defparam \always0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N30
cycloneive_lcell_comb \always0~20 (
// Equation(s):
// \always0~20_combout  = (\always0~19_combout  & (\always0~14_combout  & ((!\ramWEN~0_combout ) # (!\ramREN~0_combout ))))

	.dataa(\ramif.ramREN ),
	.datab(ramWEN),
	.datac(\always0~19_combout ),
	.datad(\always0~14_combout ),
	.cin(gnd),
	.combout(\always0~20_combout ),
	.cout());
// synopsys translate_off
defparam \always0~20 .lut_mask = 16'h7000;
defparam \always0~20 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module altsyncram_1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



altsyncram_99f1 auto_generated(
	.ram_block3a32(ram_block3a32),
	.ram_block3a0(ram_block3a0),
	.ram_block3a33(ram_block3a33),
	.ram_block3a1(ram_block3a1),
	.ram_block3a34(ram_block3a34),
	.ram_block3a2(ram_block3a2),
	.ram_block3a35(ram_block3a35),
	.ram_block3a3(ram_block3a3),
	.ram_block3a36(ram_block3a36),
	.ram_block3a4(ram_block3a4),
	.ram_block3a37(ram_block3a37),
	.ram_block3a5(ram_block3a5),
	.ram_block3a38(ram_block3a38),
	.ram_block3a6(ram_block3a6),
	.ram_block3a39(ram_block3a39),
	.ram_block3a7(ram_block3a7),
	.ram_block3a40(ram_block3a40),
	.ram_block3a8(ram_block3a8),
	.ram_block3a41(ram_block3a41),
	.ram_block3a9(ram_block3a9),
	.ram_block3a42(ram_block3a42),
	.ram_block3a10(ram_block3a10),
	.ram_block3a43(ram_block3a43),
	.ram_block3a11(ram_block3a11),
	.ram_block3a44(ram_block3a44),
	.ram_block3a12(ram_block3a12),
	.ram_block3a45(ram_block3a45),
	.ram_block3a13(ram_block3a13),
	.ram_block3a46(ram_block3a46),
	.ram_block3a14(ram_block3a14),
	.ram_block3a47(ram_block3a47),
	.ram_block3a15(ram_block3a15),
	.ram_block3a48(ram_block3a48),
	.ram_block3a16(ram_block3a16),
	.ram_block3a49(ram_block3a49),
	.ram_block3a17(ram_block3a17),
	.ram_block3a50(ram_block3a50),
	.ram_block3a18(ram_block3a18),
	.ram_block3a51(ram_block3a51),
	.ram_block3a19(ram_block3a19),
	.ram_block3a52(ram_block3a52),
	.ram_block3a20(ram_block3a20),
	.ram_block3a53(ram_block3a53),
	.ram_block3a21(ram_block3a21),
	.ram_block3a54(ram_block3a54),
	.ram_block3a22(ram_block3a22),
	.ram_block3a55(ram_block3a55),
	.ram_block3a23(ram_block3a23),
	.ram_block3a56(ram_block3a56),
	.ram_block3a24(ram_block3a24),
	.ram_block3a57(ram_block3a57),
	.ram_block3a25(ram_block3a25),
	.ram_block3a58(ram_block3a58),
	.ram_block3a26(ram_block3a26),
	.ram_block3a59(ram_block3a59),
	.ram_block3a27(ram_block3a27),
	.ram_block3a60(ram_block3a60),
	.ram_block3a28(ram_block3a28),
	.ram_block3a61(ram_block3a61),
	.ram_block3a29(ram_block3a29),
	.ram_block3a62(ram_block3a62),
	.ram_block3a30(ram_block3a30),
	.ram_block3a63(ram_block3a63),
	.ram_block3a31(ram_block3a31),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.ramaddr1(ramaddr1),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_99f1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram1|ram_block3a32~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a0~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a33~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a1~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a34~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a2~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a35~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a3~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a36~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a4~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a37~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a5~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a38~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a6~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a39~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a7~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a40~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a8~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a41~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a9~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a42~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a10~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a43~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a11~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a44~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a12~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a45~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a13~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a46~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a14~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a47~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a15~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a48~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a16~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a49~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a17~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a50~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a18~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a51~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a19~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a52~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a20~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a53~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a21~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a54~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a22~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a55~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a23~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a56~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a24~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a57~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a25~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a58~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a26~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a59~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a27~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a60~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a28~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a61~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a29~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a62~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a30~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a63~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a31~PORTBDATAOUT0 ;
wire \mgl_prim2|sdr~0_combout ;
wire [0:0] \altsyncram1|address_reg_b ;
wire [31:0] \mgl_prim2|ram_rom_data_reg ;
wire [13:0] \mgl_prim2|ram_rom_addr_reg ;


sld_mod_ram_rom mgl_prim2(
	.ram_block3a32(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a0(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a33(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a1(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a34(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a2(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a35(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a3(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a36(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a4(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a37(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a5(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a38(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a6(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a39(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a7(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a40(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a8(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a41(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a9(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a42(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a10(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a43(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a11(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a44(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a12(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a45(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a13(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a46(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a14(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a47(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a15(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a48(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a16(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a49(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a17(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a50(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a18(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a51(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a19(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a52(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a20(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a53(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a21(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a54(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a22(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a55(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a23(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a56(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a24(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a57(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a25(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a58(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a26(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a59(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a27(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a60(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a28(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a61(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a29(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a62(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a30(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a63(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a31(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.is_in_use_reg1(is_in_use_reg),
	.ram_rom_data_reg_0(\mgl_prim2|ram_rom_data_reg [0]),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.ram_rom_addr_reg_0(\mgl_prim2|ram_rom_addr_reg [0]),
	.ram_rom_addr_reg_1(\mgl_prim2|ram_rom_addr_reg [1]),
	.ram_rom_addr_reg_2(\mgl_prim2|ram_rom_addr_reg [2]),
	.ram_rom_addr_reg_3(\mgl_prim2|ram_rom_addr_reg [3]),
	.ram_rom_addr_reg_4(\mgl_prim2|ram_rom_addr_reg [4]),
	.ram_rom_addr_reg_5(\mgl_prim2|ram_rom_addr_reg [5]),
	.ram_rom_addr_reg_6(\mgl_prim2|ram_rom_addr_reg [6]),
	.ram_rom_addr_reg_7(\mgl_prim2|ram_rom_addr_reg [7]),
	.ram_rom_addr_reg_8(\mgl_prim2|ram_rom_addr_reg [8]),
	.ram_rom_addr_reg_9(\mgl_prim2|ram_rom_addr_reg [9]),
	.ram_rom_addr_reg_10(\mgl_prim2|ram_rom_addr_reg [10]),
	.ram_rom_addr_reg_11(\mgl_prim2|ram_rom_addr_reg [11]),
	.ram_rom_addr_reg_12(\mgl_prim2|ram_rom_addr_reg [12]),
	.ram_rom_data_reg_1(\mgl_prim2|ram_rom_data_reg [1]),
	.ram_rom_data_reg_2(\mgl_prim2|ram_rom_data_reg [2]),
	.ram_rom_data_reg_3(\mgl_prim2|ram_rom_data_reg [3]),
	.ram_rom_data_reg_4(\mgl_prim2|ram_rom_data_reg [4]),
	.ram_rom_data_reg_5(\mgl_prim2|ram_rom_data_reg [5]),
	.ram_rom_data_reg_6(\mgl_prim2|ram_rom_data_reg [6]),
	.ram_rom_data_reg_7(\mgl_prim2|ram_rom_data_reg [7]),
	.ram_rom_data_reg_8(\mgl_prim2|ram_rom_data_reg [8]),
	.ram_rom_data_reg_9(\mgl_prim2|ram_rom_data_reg [9]),
	.ram_rom_data_reg_10(\mgl_prim2|ram_rom_data_reg [10]),
	.ram_rom_data_reg_11(\mgl_prim2|ram_rom_data_reg [11]),
	.ram_rom_data_reg_12(\mgl_prim2|ram_rom_data_reg [12]),
	.ram_rom_data_reg_13(\mgl_prim2|ram_rom_data_reg [13]),
	.ram_rom_data_reg_14(\mgl_prim2|ram_rom_data_reg [14]),
	.ram_rom_data_reg_15(\mgl_prim2|ram_rom_data_reg [15]),
	.ram_rom_data_reg_16(\mgl_prim2|ram_rom_data_reg [16]),
	.ram_rom_data_reg_17(\mgl_prim2|ram_rom_data_reg [17]),
	.ram_rom_data_reg_18(\mgl_prim2|ram_rom_data_reg [18]),
	.ram_rom_data_reg_19(\mgl_prim2|ram_rom_data_reg [19]),
	.ram_rom_data_reg_20(\mgl_prim2|ram_rom_data_reg [20]),
	.ram_rom_data_reg_21(\mgl_prim2|ram_rom_data_reg [21]),
	.ram_rom_data_reg_22(\mgl_prim2|ram_rom_data_reg [22]),
	.ram_rom_data_reg_23(\mgl_prim2|ram_rom_data_reg [23]),
	.ram_rom_data_reg_24(\mgl_prim2|ram_rom_data_reg [24]),
	.ram_rom_data_reg_25(\mgl_prim2|ram_rom_data_reg [25]),
	.ram_rom_data_reg_26(\mgl_prim2|ram_rom_data_reg [26]),
	.ram_rom_data_reg_27(\mgl_prim2|ram_rom_data_reg [27]),
	.ram_rom_data_reg_28(\mgl_prim2|ram_rom_data_reg [28]),
	.ram_rom_data_reg_29(\mgl_prim2|ram_rom_data_reg [29]),
	.ram_rom_data_reg_30(\mgl_prim2|ram_rom_data_reg [30]),
	.ram_rom_data_reg_31(\mgl_prim2|ram_rom_data_reg [31]),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.ir_in({gnd,irf_reg_3_1,gnd,gnd,irf_reg_0_1}),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.raw_tck(altera_internal_jtag1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

altsyncram_fta2 altsyncram1(
	.ram_block3a321(ram_block3a32),
	.ram_block3a322(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a01(ram_block3a0),
	.ram_block3a02(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a331(ram_block3a33),
	.ram_block3a332(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a110(ram_block3a1),
	.ram_block3a111(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a341(ram_block3a34),
	.ram_block3a342(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a210(ram_block3a2),
	.ram_block3a211(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a351(ram_block3a35),
	.ram_block3a352(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a310(ram_block3a3),
	.ram_block3a311(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a361(ram_block3a36),
	.ram_block3a362(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a410(ram_block3a4),
	.ram_block3a411(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a371(ram_block3a37),
	.ram_block3a372(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a510(ram_block3a5),
	.ram_block3a511(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a381(ram_block3a38),
	.ram_block3a382(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a64(ram_block3a6),
	.ram_block3a65(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a391(ram_block3a39),
	.ram_block3a392(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a71(ram_block3a7),
	.ram_block3a72(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a401(ram_block3a40),
	.ram_block3a402(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a81(ram_block3a8),
	.ram_block3a82(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a412(ram_block3a41),
	.ram_block3a413(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a91(ram_block3a9),
	.ram_block3a92(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a421(ram_block3a42),
	.ram_block3a422(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a101(ram_block3a10),
	.ram_block3a102(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a431(ram_block3a43),
	.ram_block3a432(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a112(ram_block3a11),
	.ram_block3a113(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a441(ram_block3a44),
	.ram_block3a442(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a121(ram_block3a12),
	.ram_block3a122(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a451(ram_block3a45),
	.ram_block3a452(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a131(ram_block3a13),
	.ram_block3a132(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a461(ram_block3a46),
	.ram_block3a462(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a141(ram_block3a14),
	.ram_block3a142(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a471(ram_block3a47),
	.ram_block3a472(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a151(ram_block3a15),
	.ram_block3a152(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a481(ram_block3a48),
	.ram_block3a482(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a161(ram_block3a16),
	.ram_block3a162(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a491(ram_block3a49),
	.ram_block3a492(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a171(ram_block3a17),
	.ram_block3a172(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a501(ram_block3a50),
	.ram_block3a502(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a181(ram_block3a18),
	.ram_block3a182(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a512(ram_block3a51),
	.ram_block3a513(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a191(ram_block3a19),
	.ram_block3a192(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a521(ram_block3a52),
	.ram_block3a522(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a201(ram_block3a20),
	.ram_block3a202(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a531(ram_block3a53),
	.ram_block3a532(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a212(ram_block3a21),
	.ram_block3a213(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a541(ram_block3a54),
	.ram_block3a542(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a221(ram_block3a22),
	.ram_block3a222(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a551(ram_block3a55),
	.ram_block3a552(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a231(ram_block3a23),
	.ram_block3a232(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a561(ram_block3a56),
	.ram_block3a562(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a241(ram_block3a24),
	.ram_block3a242(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a571(ram_block3a57),
	.ram_block3a572(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a251(ram_block3a25),
	.ram_block3a252(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a581(ram_block3a58),
	.ram_block3a582(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a261(ram_block3a26),
	.ram_block3a262(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a591(ram_block3a59),
	.ram_block3a592(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a271(ram_block3a27),
	.ram_block3a272(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a601(ram_block3a60),
	.ram_block3a602(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a281(ram_block3a28),
	.ram_block3a282(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a611(ram_block3a61),
	.ram_block3a612(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a291(ram_block3a29),
	.ram_block3a292(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a621(ram_block3a62),
	.ram_block3a622(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a301(ram_block3a30),
	.ram_block3a302(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a631(ram_block3a63),
	.ram_block3a632(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a312(ram_block3a31),
	.ram_block3a313(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.data_b({\mgl_prim2|ram_rom_data_reg [31],\mgl_prim2|ram_rom_data_reg [30],\mgl_prim2|ram_rom_data_reg [29],\mgl_prim2|ram_rom_data_reg [28],\mgl_prim2|ram_rom_data_reg [27],\mgl_prim2|ram_rom_data_reg [26],\mgl_prim2|ram_rom_data_reg [25],\mgl_prim2|ram_rom_data_reg [24],\mgl_prim2|ram_rom_data_reg [23],
\mgl_prim2|ram_rom_data_reg [22],\mgl_prim2|ram_rom_data_reg [21],\mgl_prim2|ram_rom_data_reg [20],\mgl_prim2|ram_rom_data_reg [19],\mgl_prim2|ram_rom_data_reg [18],\mgl_prim2|ram_rom_data_reg [17],\mgl_prim2|ram_rom_data_reg [16],\mgl_prim2|ram_rom_data_reg [15],\mgl_prim2|ram_rom_data_reg [14],
\mgl_prim2|ram_rom_data_reg [13],\mgl_prim2|ram_rom_data_reg [12],\mgl_prim2|ram_rom_data_reg [11],\mgl_prim2|ram_rom_data_reg [10],\mgl_prim2|ram_rom_data_reg [9],\mgl_prim2|ram_rom_data_reg [8],\mgl_prim2|ram_rom_data_reg [7],\mgl_prim2|ram_rom_data_reg [6],\mgl_prim2|ram_rom_data_reg [5],
\mgl_prim2|ram_rom_data_reg [4],\mgl_prim2|ram_rom_data_reg [3],\mgl_prim2|ram_rom_data_reg [2],\mgl_prim2|ram_rom_data_reg [1],\mgl_prim2|ram_rom_data_reg [0]}),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.address_b({gnd,\mgl_prim2|ram_rom_addr_reg [12],\mgl_prim2|ram_rom_addr_reg [11],\mgl_prim2|ram_rom_addr_reg [10],\mgl_prim2|ram_rom_addr_reg [9],\mgl_prim2|ram_rom_addr_reg [8],\mgl_prim2|ram_rom_addr_reg [7],\mgl_prim2|ram_rom_addr_reg [6],\mgl_prim2|ram_rom_addr_reg [5],\mgl_prim2|ram_rom_addr_reg [4],
\mgl_prim2|ram_rom_addr_reg [3],\mgl_prim2|ram_rom_addr_reg [2],\mgl_prim2|ram_rom_addr_reg [1],\mgl_prim2|ram_rom_addr_reg [0]}),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.ramaddr1(ramaddr1),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.clock1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_fta2 (
	ram_block3a321,
	ram_block3a322,
	ram_block3a01,
	ram_block3a02,
	ram_block3a331,
	ram_block3a332,
	ram_block3a110,
	ram_block3a111,
	ram_block3a341,
	ram_block3a342,
	ram_block3a210,
	ram_block3a211,
	ram_block3a351,
	ram_block3a352,
	ram_block3a310,
	ram_block3a311,
	ram_block3a361,
	ram_block3a362,
	ram_block3a410,
	ram_block3a411,
	ram_block3a371,
	ram_block3a372,
	ram_block3a510,
	ram_block3a511,
	ram_block3a381,
	ram_block3a382,
	ram_block3a64,
	ram_block3a65,
	ram_block3a391,
	ram_block3a392,
	ram_block3a71,
	ram_block3a72,
	ram_block3a401,
	ram_block3a402,
	ram_block3a81,
	ram_block3a82,
	ram_block3a412,
	ram_block3a413,
	ram_block3a91,
	ram_block3a92,
	ram_block3a421,
	ram_block3a422,
	ram_block3a101,
	ram_block3a102,
	ram_block3a431,
	ram_block3a432,
	ram_block3a112,
	ram_block3a113,
	ram_block3a441,
	ram_block3a442,
	ram_block3a121,
	ram_block3a122,
	ram_block3a451,
	ram_block3a452,
	ram_block3a131,
	ram_block3a132,
	ram_block3a461,
	ram_block3a462,
	ram_block3a141,
	ram_block3a142,
	ram_block3a471,
	ram_block3a472,
	ram_block3a151,
	ram_block3a152,
	ram_block3a481,
	ram_block3a482,
	ram_block3a161,
	ram_block3a162,
	ram_block3a491,
	ram_block3a492,
	ram_block3a171,
	ram_block3a172,
	ram_block3a501,
	ram_block3a502,
	ram_block3a181,
	ram_block3a182,
	ram_block3a512,
	ram_block3a513,
	ram_block3a191,
	ram_block3a192,
	ram_block3a521,
	ram_block3a522,
	ram_block3a201,
	ram_block3a202,
	ram_block3a531,
	ram_block3a532,
	ram_block3a212,
	ram_block3a213,
	ram_block3a541,
	ram_block3a542,
	ram_block3a221,
	ram_block3a222,
	ram_block3a551,
	ram_block3a552,
	ram_block3a231,
	ram_block3a232,
	ram_block3a561,
	ram_block3a562,
	ram_block3a241,
	ram_block3a242,
	ram_block3a571,
	ram_block3a572,
	ram_block3a251,
	ram_block3a252,
	ram_block3a581,
	ram_block3a582,
	ram_block3a261,
	ram_block3a262,
	ram_block3a591,
	ram_block3a592,
	ram_block3a271,
	ram_block3a272,
	ram_block3a601,
	ram_block3a602,
	ram_block3a281,
	ram_block3a282,
	ram_block3a611,
	ram_block3a612,
	ram_block3a291,
	ram_block3a292,
	ram_block3a621,
	ram_block3a622,
	ram_block3a301,
	ram_block3a302,
	ram_block3a631,
	ram_block3a632,
	ram_block3a312,
	ram_block3a313,
	data_b,
	ram_rom_addr_reg_13,
	address_b,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	sdr,
	data_a,
	address_reg_b_0,
	ramaddr1,
	irf_reg_2_1,
	state_5,
	clock1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a321;
output 	ram_block3a322;
output 	ram_block3a01;
output 	ram_block3a02;
output 	ram_block3a331;
output 	ram_block3a332;
output 	ram_block3a110;
output 	ram_block3a111;
output 	ram_block3a341;
output 	ram_block3a342;
output 	ram_block3a210;
output 	ram_block3a211;
output 	ram_block3a351;
output 	ram_block3a352;
output 	ram_block3a310;
output 	ram_block3a311;
output 	ram_block3a361;
output 	ram_block3a362;
output 	ram_block3a410;
output 	ram_block3a411;
output 	ram_block3a371;
output 	ram_block3a372;
output 	ram_block3a510;
output 	ram_block3a511;
output 	ram_block3a381;
output 	ram_block3a382;
output 	ram_block3a64;
output 	ram_block3a65;
output 	ram_block3a391;
output 	ram_block3a392;
output 	ram_block3a71;
output 	ram_block3a72;
output 	ram_block3a401;
output 	ram_block3a402;
output 	ram_block3a81;
output 	ram_block3a82;
output 	ram_block3a412;
output 	ram_block3a413;
output 	ram_block3a91;
output 	ram_block3a92;
output 	ram_block3a421;
output 	ram_block3a422;
output 	ram_block3a101;
output 	ram_block3a102;
output 	ram_block3a431;
output 	ram_block3a432;
output 	ram_block3a112;
output 	ram_block3a113;
output 	ram_block3a441;
output 	ram_block3a442;
output 	ram_block3a121;
output 	ram_block3a122;
output 	ram_block3a451;
output 	ram_block3a452;
output 	ram_block3a131;
output 	ram_block3a132;
output 	ram_block3a461;
output 	ram_block3a462;
output 	ram_block3a141;
output 	ram_block3a142;
output 	ram_block3a471;
output 	ram_block3a472;
output 	ram_block3a151;
output 	ram_block3a152;
output 	ram_block3a481;
output 	ram_block3a482;
output 	ram_block3a161;
output 	ram_block3a162;
output 	ram_block3a491;
output 	ram_block3a492;
output 	ram_block3a171;
output 	ram_block3a172;
output 	ram_block3a501;
output 	ram_block3a502;
output 	ram_block3a181;
output 	ram_block3a182;
output 	ram_block3a512;
output 	ram_block3a513;
output 	ram_block3a191;
output 	ram_block3a192;
output 	ram_block3a521;
output 	ram_block3a522;
output 	ram_block3a201;
output 	ram_block3a202;
output 	ram_block3a531;
output 	ram_block3a532;
output 	ram_block3a212;
output 	ram_block3a213;
output 	ram_block3a541;
output 	ram_block3a542;
output 	ram_block3a221;
output 	ram_block3a222;
output 	ram_block3a551;
output 	ram_block3a552;
output 	ram_block3a231;
output 	ram_block3a232;
output 	ram_block3a561;
output 	ram_block3a562;
output 	ram_block3a241;
output 	ram_block3a242;
output 	ram_block3a571;
output 	ram_block3a572;
output 	ram_block3a251;
output 	ram_block3a252;
output 	ram_block3a581;
output 	ram_block3a582;
output 	ram_block3a261;
output 	ram_block3a262;
output 	ram_block3a591;
output 	ram_block3a592;
output 	ram_block3a271;
output 	ram_block3a272;
output 	ram_block3a601;
output 	ram_block3a602;
output 	ram_block3a281;
output 	ram_block3a282;
output 	ram_block3a611;
output 	ram_block3a612;
output 	ram_block3a291;
output 	ram_block3a292;
output 	ram_block3a621;
output 	ram_block3a622;
output 	ram_block3a301;
output 	ram_block3a302;
output 	ram_block3a631;
output 	ram_block3a632;
output 	ram_block3a312;
output 	ram_block3a313;
input 	[31:0] data_b;
input 	ram_rom_addr_reg_13;
input 	[13:0] address_b;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
input 	sdr;
input 	[31:0] data_a;
output 	address_reg_b_0;
input 	ramaddr1;
input 	irf_reg_2_1;
input 	state_5;
input 	clock1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \decode4|eq_node[1]~0_combout ;
wire \decode5|eq_node[1]~0_combout ;
wire \decode4|eq_node[0]~1_combout ;
wire \decode5|eq_node[0]~1_combout ;
wire \address_reg_b[0]~feeder_combout ;

wire [0:0] ram_block3a32_PORTADATAOUT_bus;
wire [0:0] ram_block3a32_PORTBDATAOUT_bus;
wire [0:0] ram_block3a0_PORTADATAOUT_bus;
wire [0:0] ram_block3a0_PORTBDATAOUT_bus;
wire [0:0] ram_block3a33_PORTADATAOUT_bus;
wire [0:0] ram_block3a33_PORTBDATAOUT_bus;
wire [0:0] ram_block3a1_PORTADATAOUT_bus;
wire [0:0] ram_block3a1_PORTBDATAOUT_bus;
wire [0:0] ram_block3a34_PORTADATAOUT_bus;
wire [0:0] ram_block3a34_PORTBDATAOUT_bus;
wire [0:0] ram_block3a2_PORTADATAOUT_bus;
wire [0:0] ram_block3a2_PORTBDATAOUT_bus;
wire [0:0] ram_block3a35_PORTADATAOUT_bus;
wire [0:0] ram_block3a35_PORTBDATAOUT_bus;
wire [0:0] ram_block3a3_PORTADATAOUT_bus;
wire [0:0] ram_block3a3_PORTBDATAOUT_bus;
wire [0:0] ram_block3a36_PORTADATAOUT_bus;
wire [0:0] ram_block3a36_PORTBDATAOUT_bus;
wire [0:0] ram_block3a4_PORTADATAOUT_bus;
wire [0:0] ram_block3a4_PORTBDATAOUT_bus;
wire [0:0] ram_block3a37_PORTADATAOUT_bus;
wire [0:0] ram_block3a37_PORTBDATAOUT_bus;
wire [0:0] ram_block3a5_PORTADATAOUT_bus;
wire [0:0] ram_block3a5_PORTBDATAOUT_bus;
wire [0:0] ram_block3a38_PORTADATAOUT_bus;
wire [0:0] ram_block3a38_PORTBDATAOUT_bus;
wire [0:0] ram_block3a6_PORTADATAOUT_bus;
wire [0:0] ram_block3a6_PORTBDATAOUT_bus;
wire [0:0] ram_block3a39_PORTADATAOUT_bus;
wire [0:0] ram_block3a39_PORTBDATAOUT_bus;
wire [0:0] ram_block3a7_PORTADATAOUT_bus;
wire [0:0] ram_block3a7_PORTBDATAOUT_bus;
wire [0:0] ram_block3a40_PORTADATAOUT_bus;
wire [0:0] ram_block3a40_PORTBDATAOUT_bus;
wire [0:0] ram_block3a8_PORTADATAOUT_bus;
wire [0:0] ram_block3a8_PORTBDATAOUT_bus;
wire [0:0] ram_block3a41_PORTADATAOUT_bus;
wire [0:0] ram_block3a41_PORTBDATAOUT_bus;
wire [0:0] ram_block3a9_PORTADATAOUT_bus;
wire [0:0] ram_block3a9_PORTBDATAOUT_bus;
wire [0:0] ram_block3a42_PORTADATAOUT_bus;
wire [0:0] ram_block3a42_PORTBDATAOUT_bus;
wire [0:0] ram_block3a10_PORTADATAOUT_bus;
wire [0:0] ram_block3a10_PORTBDATAOUT_bus;
wire [0:0] ram_block3a43_PORTADATAOUT_bus;
wire [0:0] ram_block3a43_PORTBDATAOUT_bus;
wire [0:0] ram_block3a11_PORTADATAOUT_bus;
wire [0:0] ram_block3a11_PORTBDATAOUT_bus;
wire [0:0] ram_block3a44_PORTADATAOUT_bus;
wire [0:0] ram_block3a44_PORTBDATAOUT_bus;
wire [0:0] ram_block3a12_PORTADATAOUT_bus;
wire [0:0] ram_block3a12_PORTBDATAOUT_bus;
wire [0:0] ram_block3a45_PORTADATAOUT_bus;
wire [0:0] ram_block3a45_PORTBDATAOUT_bus;
wire [0:0] ram_block3a13_PORTADATAOUT_bus;
wire [0:0] ram_block3a13_PORTBDATAOUT_bus;
wire [0:0] ram_block3a46_PORTADATAOUT_bus;
wire [0:0] ram_block3a46_PORTBDATAOUT_bus;
wire [0:0] ram_block3a14_PORTADATAOUT_bus;
wire [0:0] ram_block3a14_PORTBDATAOUT_bus;
wire [0:0] ram_block3a47_PORTADATAOUT_bus;
wire [0:0] ram_block3a47_PORTBDATAOUT_bus;
wire [0:0] ram_block3a15_PORTADATAOUT_bus;
wire [0:0] ram_block3a15_PORTBDATAOUT_bus;
wire [0:0] ram_block3a48_PORTADATAOUT_bus;
wire [0:0] ram_block3a48_PORTBDATAOUT_bus;
wire [0:0] ram_block3a16_PORTADATAOUT_bus;
wire [0:0] ram_block3a16_PORTBDATAOUT_bus;
wire [0:0] ram_block3a49_PORTADATAOUT_bus;
wire [0:0] ram_block3a49_PORTBDATAOUT_bus;
wire [0:0] ram_block3a17_PORTADATAOUT_bus;
wire [0:0] ram_block3a17_PORTBDATAOUT_bus;
wire [0:0] ram_block3a50_PORTADATAOUT_bus;
wire [0:0] ram_block3a50_PORTBDATAOUT_bus;
wire [0:0] ram_block3a18_PORTADATAOUT_bus;
wire [0:0] ram_block3a18_PORTBDATAOUT_bus;
wire [0:0] ram_block3a51_PORTADATAOUT_bus;
wire [0:0] ram_block3a51_PORTBDATAOUT_bus;
wire [0:0] ram_block3a19_PORTADATAOUT_bus;
wire [0:0] ram_block3a19_PORTBDATAOUT_bus;
wire [0:0] ram_block3a52_PORTADATAOUT_bus;
wire [0:0] ram_block3a52_PORTBDATAOUT_bus;
wire [0:0] ram_block3a20_PORTADATAOUT_bus;
wire [0:0] ram_block3a20_PORTBDATAOUT_bus;
wire [0:0] ram_block3a53_PORTADATAOUT_bus;
wire [0:0] ram_block3a53_PORTBDATAOUT_bus;
wire [0:0] ram_block3a21_PORTADATAOUT_bus;
wire [0:0] ram_block3a21_PORTBDATAOUT_bus;
wire [0:0] ram_block3a54_PORTADATAOUT_bus;
wire [0:0] ram_block3a54_PORTBDATAOUT_bus;
wire [0:0] ram_block3a22_PORTADATAOUT_bus;
wire [0:0] ram_block3a22_PORTBDATAOUT_bus;
wire [0:0] ram_block3a55_PORTADATAOUT_bus;
wire [0:0] ram_block3a55_PORTBDATAOUT_bus;
wire [0:0] ram_block3a23_PORTADATAOUT_bus;
wire [0:0] ram_block3a23_PORTBDATAOUT_bus;
wire [0:0] ram_block3a56_PORTADATAOUT_bus;
wire [0:0] ram_block3a56_PORTBDATAOUT_bus;
wire [0:0] ram_block3a24_PORTADATAOUT_bus;
wire [0:0] ram_block3a24_PORTBDATAOUT_bus;
wire [0:0] ram_block3a57_PORTADATAOUT_bus;
wire [0:0] ram_block3a57_PORTBDATAOUT_bus;
wire [0:0] ram_block3a25_PORTADATAOUT_bus;
wire [0:0] ram_block3a25_PORTBDATAOUT_bus;
wire [0:0] ram_block3a58_PORTADATAOUT_bus;
wire [0:0] ram_block3a58_PORTBDATAOUT_bus;
wire [0:0] ram_block3a26_PORTADATAOUT_bus;
wire [0:0] ram_block3a26_PORTBDATAOUT_bus;
wire [0:0] ram_block3a59_PORTADATAOUT_bus;
wire [0:0] ram_block3a59_PORTBDATAOUT_bus;
wire [0:0] ram_block3a27_PORTADATAOUT_bus;
wire [0:0] ram_block3a27_PORTBDATAOUT_bus;
wire [0:0] ram_block3a60_PORTADATAOUT_bus;
wire [0:0] ram_block3a60_PORTBDATAOUT_bus;
wire [0:0] ram_block3a28_PORTADATAOUT_bus;
wire [0:0] ram_block3a28_PORTBDATAOUT_bus;
wire [0:0] ram_block3a61_PORTADATAOUT_bus;
wire [0:0] ram_block3a61_PORTBDATAOUT_bus;
wire [0:0] ram_block3a29_PORTADATAOUT_bus;
wire [0:0] ram_block3a29_PORTBDATAOUT_bus;
wire [0:0] ram_block3a62_PORTADATAOUT_bus;
wire [0:0] ram_block3a62_PORTBDATAOUT_bus;
wire [0:0] ram_block3a30_PORTADATAOUT_bus;
wire [0:0] ram_block3a30_PORTBDATAOUT_bus;
wire [0:0] ram_block3a63_PORTADATAOUT_bus;
wire [0:0] ram_block3a63_PORTBDATAOUT_bus;
wire [0:0] ram_block3a31_PORTADATAOUT_bus;
wire [0:0] ram_block3a31_PORTBDATAOUT_bus;

assign ram_block3a321 = ram_block3a32_PORTADATAOUT_bus[0];

assign ram_block3a322 = ram_block3a32_PORTBDATAOUT_bus[0];

assign ram_block3a01 = ram_block3a0_PORTADATAOUT_bus[0];

assign ram_block3a02 = ram_block3a0_PORTBDATAOUT_bus[0];

assign ram_block3a331 = ram_block3a33_PORTADATAOUT_bus[0];

assign ram_block3a332 = ram_block3a33_PORTBDATAOUT_bus[0];

assign ram_block3a110 = ram_block3a1_PORTADATAOUT_bus[0];

assign ram_block3a111 = ram_block3a1_PORTBDATAOUT_bus[0];

assign ram_block3a341 = ram_block3a34_PORTADATAOUT_bus[0];

assign ram_block3a342 = ram_block3a34_PORTBDATAOUT_bus[0];

assign ram_block3a210 = ram_block3a2_PORTADATAOUT_bus[0];

assign ram_block3a211 = ram_block3a2_PORTBDATAOUT_bus[0];

assign ram_block3a351 = ram_block3a35_PORTADATAOUT_bus[0];

assign ram_block3a352 = ram_block3a35_PORTBDATAOUT_bus[0];

assign ram_block3a310 = ram_block3a3_PORTADATAOUT_bus[0];

assign ram_block3a311 = ram_block3a3_PORTBDATAOUT_bus[0];

assign ram_block3a361 = ram_block3a36_PORTADATAOUT_bus[0];

assign ram_block3a362 = ram_block3a36_PORTBDATAOUT_bus[0];

assign ram_block3a410 = ram_block3a4_PORTADATAOUT_bus[0];

assign ram_block3a411 = ram_block3a4_PORTBDATAOUT_bus[0];

assign ram_block3a371 = ram_block3a37_PORTADATAOUT_bus[0];

assign ram_block3a372 = ram_block3a37_PORTBDATAOUT_bus[0];

assign ram_block3a510 = ram_block3a5_PORTADATAOUT_bus[0];

assign ram_block3a511 = ram_block3a5_PORTBDATAOUT_bus[0];

assign ram_block3a381 = ram_block3a38_PORTADATAOUT_bus[0];

assign ram_block3a382 = ram_block3a38_PORTBDATAOUT_bus[0];

assign ram_block3a64 = ram_block3a6_PORTADATAOUT_bus[0];

assign ram_block3a65 = ram_block3a6_PORTBDATAOUT_bus[0];

assign ram_block3a391 = ram_block3a39_PORTADATAOUT_bus[0];

assign ram_block3a392 = ram_block3a39_PORTBDATAOUT_bus[0];

assign ram_block3a71 = ram_block3a7_PORTADATAOUT_bus[0];

assign ram_block3a72 = ram_block3a7_PORTBDATAOUT_bus[0];

assign ram_block3a401 = ram_block3a40_PORTADATAOUT_bus[0];

assign ram_block3a402 = ram_block3a40_PORTBDATAOUT_bus[0];

assign ram_block3a81 = ram_block3a8_PORTADATAOUT_bus[0];

assign ram_block3a82 = ram_block3a8_PORTBDATAOUT_bus[0];

assign ram_block3a412 = ram_block3a41_PORTADATAOUT_bus[0];

assign ram_block3a413 = ram_block3a41_PORTBDATAOUT_bus[0];

assign ram_block3a91 = ram_block3a9_PORTADATAOUT_bus[0];

assign ram_block3a92 = ram_block3a9_PORTBDATAOUT_bus[0];

assign ram_block3a421 = ram_block3a42_PORTADATAOUT_bus[0];

assign ram_block3a422 = ram_block3a42_PORTBDATAOUT_bus[0];

assign ram_block3a101 = ram_block3a10_PORTADATAOUT_bus[0];

assign ram_block3a102 = ram_block3a10_PORTBDATAOUT_bus[0];

assign ram_block3a431 = ram_block3a43_PORTADATAOUT_bus[0];

assign ram_block3a432 = ram_block3a43_PORTBDATAOUT_bus[0];

assign ram_block3a112 = ram_block3a11_PORTADATAOUT_bus[0];

assign ram_block3a113 = ram_block3a11_PORTBDATAOUT_bus[0];

assign ram_block3a441 = ram_block3a44_PORTADATAOUT_bus[0];

assign ram_block3a442 = ram_block3a44_PORTBDATAOUT_bus[0];

assign ram_block3a121 = ram_block3a12_PORTADATAOUT_bus[0];

assign ram_block3a122 = ram_block3a12_PORTBDATAOUT_bus[0];

assign ram_block3a451 = ram_block3a45_PORTADATAOUT_bus[0];

assign ram_block3a452 = ram_block3a45_PORTBDATAOUT_bus[0];

assign ram_block3a131 = ram_block3a13_PORTADATAOUT_bus[0];

assign ram_block3a132 = ram_block3a13_PORTBDATAOUT_bus[0];

assign ram_block3a461 = ram_block3a46_PORTADATAOUT_bus[0];

assign ram_block3a462 = ram_block3a46_PORTBDATAOUT_bus[0];

assign ram_block3a141 = ram_block3a14_PORTADATAOUT_bus[0];

assign ram_block3a142 = ram_block3a14_PORTBDATAOUT_bus[0];

assign ram_block3a471 = ram_block3a47_PORTADATAOUT_bus[0];

assign ram_block3a472 = ram_block3a47_PORTBDATAOUT_bus[0];

assign ram_block3a151 = ram_block3a15_PORTADATAOUT_bus[0];

assign ram_block3a152 = ram_block3a15_PORTBDATAOUT_bus[0];

assign ram_block3a481 = ram_block3a48_PORTADATAOUT_bus[0];

assign ram_block3a482 = ram_block3a48_PORTBDATAOUT_bus[0];

assign ram_block3a161 = ram_block3a16_PORTADATAOUT_bus[0];

assign ram_block3a162 = ram_block3a16_PORTBDATAOUT_bus[0];

assign ram_block3a491 = ram_block3a49_PORTADATAOUT_bus[0];

assign ram_block3a492 = ram_block3a49_PORTBDATAOUT_bus[0];

assign ram_block3a171 = ram_block3a17_PORTADATAOUT_bus[0];

assign ram_block3a172 = ram_block3a17_PORTBDATAOUT_bus[0];

assign ram_block3a501 = ram_block3a50_PORTADATAOUT_bus[0];

assign ram_block3a502 = ram_block3a50_PORTBDATAOUT_bus[0];

assign ram_block3a181 = ram_block3a18_PORTADATAOUT_bus[0];

assign ram_block3a182 = ram_block3a18_PORTBDATAOUT_bus[0];

assign ram_block3a512 = ram_block3a51_PORTADATAOUT_bus[0];

assign ram_block3a513 = ram_block3a51_PORTBDATAOUT_bus[0];

assign ram_block3a191 = ram_block3a19_PORTADATAOUT_bus[0];

assign ram_block3a192 = ram_block3a19_PORTBDATAOUT_bus[0];

assign ram_block3a521 = ram_block3a52_PORTADATAOUT_bus[0];

assign ram_block3a522 = ram_block3a52_PORTBDATAOUT_bus[0];

assign ram_block3a201 = ram_block3a20_PORTADATAOUT_bus[0];

assign ram_block3a202 = ram_block3a20_PORTBDATAOUT_bus[0];

assign ram_block3a531 = ram_block3a53_PORTADATAOUT_bus[0];

assign ram_block3a532 = ram_block3a53_PORTBDATAOUT_bus[0];

assign ram_block3a212 = ram_block3a21_PORTADATAOUT_bus[0];

assign ram_block3a213 = ram_block3a21_PORTBDATAOUT_bus[0];

assign ram_block3a541 = ram_block3a54_PORTADATAOUT_bus[0];

assign ram_block3a542 = ram_block3a54_PORTBDATAOUT_bus[0];

assign ram_block3a221 = ram_block3a22_PORTADATAOUT_bus[0];

assign ram_block3a222 = ram_block3a22_PORTBDATAOUT_bus[0];

assign ram_block3a551 = ram_block3a55_PORTADATAOUT_bus[0];

assign ram_block3a552 = ram_block3a55_PORTBDATAOUT_bus[0];

assign ram_block3a231 = ram_block3a23_PORTADATAOUT_bus[0];

assign ram_block3a232 = ram_block3a23_PORTBDATAOUT_bus[0];

assign ram_block3a561 = ram_block3a56_PORTADATAOUT_bus[0];

assign ram_block3a562 = ram_block3a56_PORTBDATAOUT_bus[0];

assign ram_block3a241 = ram_block3a24_PORTADATAOUT_bus[0];

assign ram_block3a242 = ram_block3a24_PORTBDATAOUT_bus[0];

assign ram_block3a571 = ram_block3a57_PORTADATAOUT_bus[0];

assign ram_block3a572 = ram_block3a57_PORTBDATAOUT_bus[0];

assign ram_block3a251 = ram_block3a25_PORTADATAOUT_bus[0];

assign ram_block3a252 = ram_block3a25_PORTBDATAOUT_bus[0];

assign ram_block3a581 = ram_block3a58_PORTADATAOUT_bus[0];

assign ram_block3a582 = ram_block3a58_PORTBDATAOUT_bus[0];

assign ram_block3a261 = ram_block3a26_PORTADATAOUT_bus[0];

assign ram_block3a262 = ram_block3a26_PORTBDATAOUT_bus[0];

assign ram_block3a591 = ram_block3a59_PORTADATAOUT_bus[0];

assign ram_block3a592 = ram_block3a59_PORTBDATAOUT_bus[0];

assign ram_block3a271 = ram_block3a27_PORTADATAOUT_bus[0];

assign ram_block3a272 = ram_block3a27_PORTBDATAOUT_bus[0];

assign ram_block3a601 = ram_block3a60_PORTADATAOUT_bus[0];

assign ram_block3a602 = ram_block3a60_PORTBDATAOUT_bus[0];

assign ram_block3a281 = ram_block3a28_PORTADATAOUT_bus[0];

assign ram_block3a282 = ram_block3a28_PORTBDATAOUT_bus[0];

assign ram_block3a611 = ram_block3a61_PORTADATAOUT_bus[0];

assign ram_block3a612 = ram_block3a61_PORTBDATAOUT_bus[0];

assign ram_block3a291 = ram_block3a29_PORTADATAOUT_bus[0];

assign ram_block3a292 = ram_block3a29_PORTBDATAOUT_bus[0];

assign ram_block3a621 = ram_block3a62_PORTADATAOUT_bus[0];

assign ram_block3a622 = ram_block3a62_PORTBDATAOUT_bus[0];

assign ram_block3a301 = ram_block3a30_PORTADATAOUT_bus[0];

assign ram_block3a302 = ram_block3a30_PORTBDATAOUT_bus[0];

assign ram_block3a631 = ram_block3a63_PORTADATAOUT_bus[0];

assign ram_block3a632 = ram_block3a63_PORTBDATAOUT_bus[0];

assign ram_block3a312 = ram_block3a31_PORTADATAOUT_bus[0];

assign ram_block3a313 = ram_block3a31_PORTBDATAOUT_bus[0];

decode_jsa_1 decode5(
	.ram_rom_addr_reg_13(ram_rom_addr_reg_13),
	.sdr(sdr),
	.eq_node_1(\decode5|eq_node[1]~0_combout ),
	.eq_node_0(\decode5|eq_node[0]~1_combout ),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

decode_jsa decode4(
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.eq_node_1(\decode4|eq_node[1]~0_combout ),
	.eq_node_0(\decode4|eq_node[0]~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: M9K_X37_Y35_N0
cycloneive_ram_block ram_block3a32(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a32_PORTADATAOUT_bus),
	.portbdataout(ram_block3a32_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a32.clk0_core_clock_enable = "ena0";
defparam ram_block3a32.clk1_core_clock_enable = "ena1";
defparam ram_block3a32.data_interleave_offset_in_bits = 1;
defparam ram_block3a32.data_interleave_width_in_bits = 1;
defparam ram_block3a32.init_file = "meminit.hex";
defparam ram_block3a32.init_file_layout = "port_a";
defparam ram_block3a32.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a32.operation_mode = "bidir_dual_port";
defparam ram_block3a32.port_a_address_clear = "none";
defparam ram_block3a32.port_a_address_width = 13;
defparam ram_block3a32.port_a_byte_enable_clock = "none";
defparam ram_block3a32.port_a_data_out_clear = "none";
defparam ram_block3a32.port_a_data_out_clock = "none";
defparam ram_block3a32.port_a_data_width = 1;
defparam ram_block3a32.port_a_first_address = 0;
defparam ram_block3a32.port_a_first_bit_number = 0;
defparam ram_block3a32.port_a_last_address = 8191;
defparam ram_block3a32.port_a_logical_ram_depth = 16384;
defparam ram_block3a32.port_a_logical_ram_width = 32;
defparam ram_block3a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_address_clear = "none";
defparam ram_block3a32.port_b_address_clock = "clock1";
defparam ram_block3a32.port_b_address_width = 13;
defparam ram_block3a32.port_b_data_in_clock = "clock1";
defparam ram_block3a32.port_b_data_out_clear = "none";
defparam ram_block3a32.port_b_data_out_clock = "none";
defparam ram_block3a32.port_b_data_width = 1;
defparam ram_block3a32.port_b_first_address = 0;
defparam ram_block3a32.port_b_first_bit_number = 0;
defparam ram_block3a32.port_b_last_address = 8191;
defparam ram_block3a32.port_b_logical_ram_depth = 16384;
defparam ram_block3a32.port_b_logical_ram_width = 32;
defparam ram_block3a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_read_enable_clock = "clock1";
defparam ram_block3a32.port_b_write_enable_clock = "clock1";
defparam ram_block3a32.ram_block_type = "M9K";
defparam ram_block3a32.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y34_N0
cycloneive_ram_block ram_block3a0(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a0_PORTADATAOUT_bus),
	.portbdataout(ram_block3a0_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a0.clk0_core_clock_enable = "ena0";
defparam ram_block3a0.clk1_core_clock_enable = "ena1";
defparam ram_block3a0.data_interleave_offset_in_bits = 1;
defparam ram_block3a0.data_interleave_width_in_bits = 1;
defparam ram_block3a0.init_file = "meminit.hex";
defparam ram_block3a0.init_file_layout = "port_a";
defparam ram_block3a0.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a0.operation_mode = "bidir_dual_port";
defparam ram_block3a0.port_a_address_clear = "none";
defparam ram_block3a0.port_a_address_width = 13;
defparam ram_block3a0.port_a_byte_enable_clock = "none";
defparam ram_block3a0.port_a_data_out_clear = "none";
defparam ram_block3a0.port_a_data_out_clock = "none";
defparam ram_block3a0.port_a_data_width = 1;
defparam ram_block3a0.port_a_first_address = 0;
defparam ram_block3a0.port_a_first_bit_number = 0;
defparam ram_block3a0.port_a_last_address = 8191;
defparam ram_block3a0.port_a_logical_ram_depth = 16384;
defparam ram_block3a0.port_a_logical_ram_width = 32;
defparam ram_block3a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_address_clear = "none";
defparam ram_block3a0.port_b_address_clock = "clock1";
defparam ram_block3a0.port_b_address_width = 13;
defparam ram_block3a0.port_b_data_in_clock = "clock1";
defparam ram_block3a0.port_b_data_out_clear = "none";
defparam ram_block3a0.port_b_data_out_clock = "none";
defparam ram_block3a0.port_b_data_width = 1;
defparam ram_block3a0.port_b_first_address = 0;
defparam ram_block3a0.port_b_first_bit_number = 0;
defparam ram_block3a0.port_b_last_address = 8191;
defparam ram_block3a0.port_b_logical_ram_depth = 16384;
defparam ram_block3a0.port_b_logical_ram_width = 32;
defparam ram_block3a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_read_enable_clock = "clock1";
defparam ram_block3a0.port_b_write_enable_clock = "clock1";
defparam ram_block3a0.ram_block_type = "M9K";
defparam ram_block3a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001802C7EA14A7EF95C00000000000000000000000000000A242111E008528F7260;
// synopsys translate_on

// Location: M9K_X64_Y39_N0
cycloneive_ram_block ram_block3a33(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a33_PORTADATAOUT_bus),
	.portbdataout(ram_block3a33_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a33.clk0_core_clock_enable = "ena0";
defparam ram_block3a33.clk1_core_clock_enable = "ena1";
defparam ram_block3a33.data_interleave_offset_in_bits = 1;
defparam ram_block3a33.data_interleave_width_in_bits = 1;
defparam ram_block3a33.init_file = "meminit.hex";
defparam ram_block3a33.init_file_layout = "port_a";
defparam ram_block3a33.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a33.operation_mode = "bidir_dual_port";
defparam ram_block3a33.port_a_address_clear = "none";
defparam ram_block3a33.port_a_address_width = 13;
defparam ram_block3a33.port_a_byte_enable_clock = "none";
defparam ram_block3a33.port_a_data_out_clear = "none";
defparam ram_block3a33.port_a_data_out_clock = "none";
defparam ram_block3a33.port_a_data_width = 1;
defparam ram_block3a33.port_a_first_address = 0;
defparam ram_block3a33.port_a_first_bit_number = 1;
defparam ram_block3a33.port_a_last_address = 8191;
defparam ram_block3a33.port_a_logical_ram_depth = 16384;
defparam ram_block3a33.port_a_logical_ram_width = 32;
defparam ram_block3a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_address_clear = "none";
defparam ram_block3a33.port_b_address_clock = "clock1";
defparam ram_block3a33.port_b_address_width = 13;
defparam ram_block3a33.port_b_data_in_clock = "clock1";
defparam ram_block3a33.port_b_data_out_clear = "none";
defparam ram_block3a33.port_b_data_out_clock = "none";
defparam ram_block3a33.port_b_data_width = 1;
defparam ram_block3a33.port_b_first_address = 0;
defparam ram_block3a33.port_b_first_bit_number = 1;
defparam ram_block3a33.port_b_last_address = 8191;
defparam ram_block3a33.port_b_logical_ram_depth = 16384;
defparam ram_block3a33.port_b_logical_ram_width = 32;
defparam ram_block3a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_read_enable_clock = "clock1";
defparam ram_block3a33.port_b_write_enable_clock = "clock1";
defparam ram_block3a33.ram_block_type = "M9K";
defparam ram_block3a33.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y38_N0
cycloneive_ram_block ram_block3a1(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a1_PORTADATAOUT_bus),
	.portbdataout(ram_block3a1_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a1.clk0_core_clock_enable = "ena0";
defparam ram_block3a1.clk1_core_clock_enable = "ena1";
defparam ram_block3a1.data_interleave_offset_in_bits = 1;
defparam ram_block3a1.data_interleave_width_in_bits = 1;
defparam ram_block3a1.init_file = "meminit.hex";
defparam ram_block3a1.init_file_layout = "port_a";
defparam ram_block3a1.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a1.operation_mode = "bidir_dual_port";
defparam ram_block3a1.port_a_address_clear = "none";
defparam ram_block3a1.port_a_address_width = 13;
defparam ram_block3a1.port_a_byte_enable_clock = "none";
defparam ram_block3a1.port_a_data_out_clear = "none";
defparam ram_block3a1.port_a_data_out_clock = "none";
defparam ram_block3a1.port_a_data_width = 1;
defparam ram_block3a1.port_a_first_address = 0;
defparam ram_block3a1.port_a_first_bit_number = 1;
defparam ram_block3a1.port_a_last_address = 8191;
defparam ram_block3a1.port_a_logical_ram_depth = 16384;
defparam ram_block3a1.port_a_logical_ram_width = 32;
defparam ram_block3a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_address_clear = "none";
defparam ram_block3a1.port_b_address_clock = "clock1";
defparam ram_block3a1.port_b_address_width = 13;
defparam ram_block3a1.port_b_data_in_clock = "clock1";
defparam ram_block3a1.port_b_data_out_clear = "none";
defparam ram_block3a1.port_b_data_out_clock = "none";
defparam ram_block3a1.port_b_data_width = 1;
defparam ram_block3a1.port_b_first_address = 0;
defparam ram_block3a1.port_b_first_bit_number = 1;
defparam ram_block3a1.port_b_last_address = 8191;
defparam ram_block3a1.port_b_logical_ram_depth = 16384;
defparam ram_block3a1.port_b_logical_ram_width = 32;
defparam ram_block3a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_read_enable_clock = "clock1";
defparam ram_block3a1.port_b_write_enable_clock = "clock1";
defparam ram_block3a1.ram_block_type = "M9K";
defparam ram_block3a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001D4AE6429116B3C8A000000000000000000000000000012242108900D12808390;
// synopsys translate_on

// Location: M9K_X64_Y40_N0
cycloneive_ram_block ram_block3a34(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a34_PORTADATAOUT_bus),
	.portbdataout(ram_block3a34_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a34.clk0_core_clock_enable = "ena0";
defparam ram_block3a34.clk1_core_clock_enable = "ena1";
defparam ram_block3a34.data_interleave_offset_in_bits = 1;
defparam ram_block3a34.data_interleave_width_in_bits = 1;
defparam ram_block3a34.init_file = "meminit.hex";
defparam ram_block3a34.init_file_layout = "port_a";
defparam ram_block3a34.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a34.operation_mode = "bidir_dual_port";
defparam ram_block3a34.port_a_address_clear = "none";
defparam ram_block3a34.port_a_address_width = 13;
defparam ram_block3a34.port_a_byte_enable_clock = "none";
defparam ram_block3a34.port_a_data_out_clear = "none";
defparam ram_block3a34.port_a_data_out_clock = "none";
defparam ram_block3a34.port_a_data_width = 1;
defparam ram_block3a34.port_a_first_address = 0;
defparam ram_block3a34.port_a_first_bit_number = 2;
defparam ram_block3a34.port_a_last_address = 8191;
defparam ram_block3a34.port_a_logical_ram_depth = 16384;
defparam ram_block3a34.port_a_logical_ram_width = 32;
defparam ram_block3a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_address_clear = "none";
defparam ram_block3a34.port_b_address_clock = "clock1";
defparam ram_block3a34.port_b_address_width = 13;
defparam ram_block3a34.port_b_data_in_clock = "clock1";
defparam ram_block3a34.port_b_data_out_clear = "none";
defparam ram_block3a34.port_b_data_out_clock = "none";
defparam ram_block3a34.port_b_data_width = 1;
defparam ram_block3a34.port_b_first_address = 0;
defparam ram_block3a34.port_b_first_bit_number = 2;
defparam ram_block3a34.port_b_last_address = 8191;
defparam ram_block3a34.port_b_logical_ram_depth = 16384;
defparam ram_block3a34.port_b_logical_ram_width = 32;
defparam ram_block3a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_read_enable_clock = "clock1";
defparam ram_block3a34.port_b_write_enable_clock = "clock1";
defparam ram_block3a34.ram_block_type = "M9K";
defparam ram_block3a34.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y41_N0
cycloneive_ram_block ram_block3a2(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a2_PORTADATAOUT_bus),
	.portbdataout(ram_block3a2_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a2.clk0_core_clock_enable = "ena0";
defparam ram_block3a2.clk1_core_clock_enable = "ena1";
defparam ram_block3a2.data_interleave_offset_in_bits = 1;
defparam ram_block3a2.data_interleave_width_in_bits = 1;
defparam ram_block3a2.init_file = "meminit.hex";
defparam ram_block3a2.init_file_layout = "port_a";
defparam ram_block3a2.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a2.operation_mode = "bidir_dual_port";
defparam ram_block3a2.port_a_address_clear = "none";
defparam ram_block3a2.port_a_address_width = 13;
defparam ram_block3a2.port_a_byte_enable_clock = "none";
defparam ram_block3a2.port_a_data_out_clear = "none";
defparam ram_block3a2.port_a_data_out_clock = "none";
defparam ram_block3a2.port_a_data_width = 1;
defparam ram_block3a2.port_a_first_address = 0;
defparam ram_block3a2.port_a_first_bit_number = 2;
defparam ram_block3a2.port_a_last_address = 8191;
defparam ram_block3a2.port_a_logical_ram_depth = 16384;
defparam ram_block3a2.port_a_logical_ram_width = 32;
defparam ram_block3a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_address_clear = "none";
defparam ram_block3a2.port_b_address_clock = "clock1";
defparam ram_block3a2.port_b_address_width = 13;
defparam ram_block3a2.port_b_data_in_clock = "clock1";
defparam ram_block3a2.port_b_data_out_clear = "none";
defparam ram_block3a2.port_b_data_out_clock = "none";
defparam ram_block3a2.port_b_data_width = 1;
defparam ram_block3a2.port_b_first_address = 0;
defparam ram_block3a2.port_b_first_bit_number = 2;
defparam ram_block3a2.port_b_last_address = 8191;
defparam ram_block3a2.port_b_logical_ram_depth = 16384;
defparam ram_block3a2.port_b_logical_ram_width = 32;
defparam ram_block3a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_read_enable_clock = "clock1";
defparam ram_block3a2.port_b_write_enable_clock = "clock1";
defparam ram_block3a2.ram_block_type = "M9K";
defparam ram_block3a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000961CA470728D97800000000000000000000000000000172E7BD1C323272F6867;
// synopsys translate_on

// Location: M9K_X37_Y36_N0
cycloneive_ram_block ram_block3a35(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a35_PORTADATAOUT_bus),
	.portbdataout(ram_block3a35_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a35.clk0_core_clock_enable = "ena0";
defparam ram_block3a35.clk1_core_clock_enable = "ena1";
defparam ram_block3a35.data_interleave_offset_in_bits = 1;
defparam ram_block3a35.data_interleave_width_in_bits = 1;
defparam ram_block3a35.init_file = "meminit.hex";
defparam ram_block3a35.init_file_layout = "port_a";
defparam ram_block3a35.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a35.operation_mode = "bidir_dual_port";
defparam ram_block3a35.port_a_address_clear = "none";
defparam ram_block3a35.port_a_address_width = 13;
defparam ram_block3a35.port_a_byte_enable_clock = "none";
defparam ram_block3a35.port_a_data_out_clear = "none";
defparam ram_block3a35.port_a_data_out_clock = "none";
defparam ram_block3a35.port_a_data_width = 1;
defparam ram_block3a35.port_a_first_address = 0;
defparam ram_block3a35.port_a_first_bit_number = 3;
defparam ram_block3a35.port_a_last_address = 8191;
defparam ram_block3a35.port_a_logical_ram_depth = 16384;
defparam ram_block3a35.port_a_logical_ram_width = 32;
defparam ram_block3a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_address_clear = "none";
defparam ram_block3a35.port_b_address_clock = "clock1";
defparam ram_block3a35.port_b_address_width = 13;
defparam ram_block3a35.port_b_data_in_clock = "clock1";
defparam ram_block3a35.port_b_data_out_clear = "none";
defparam ram_block3a35.port_b_data_out_clock = "none";
defparam ram_block3a35.port_b_data_width = 1;
defparam ram_block3a35.port_b_first_address = 0;
defparam ram_block3a35.port_b_first_bit_number = 3;
defparam ram_block3a35.port_b_last_address = 8191;
defparam ram_block3a35.port_b_logical_ram_depth = 16384;
defparam ram_block3a35.port_b_logical_ram_width = 32;
defparam ram_block3a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_read_enable_clock = "clock1";
defparam ram_block3a35.port_b_write_enable_clock = "clock1";
defparam ram_block3a35.ram_block_type = "M9K";
defparam ram_block3a35.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y36_N0
cycloneive_ram_block ram_block3a3(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a3_PORTADATAOUT_bus),
	.portbdataout(ram_block3a3_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a3.clk0_core_clock_enable = "ena0";
defparam ram_block3a3.clk1_core_clock_enable = "ena1";
defparam ram_block3a3.data_interleave_offset_in_bits = 1;
defparam ram_block3a3.data_interleave_width_in_bits = 1;
defparam ram_block3a3.init_file = "meminit.hex";
defparam ram_block3a3.init_file_layout = "port_a";
defparam ram_block3a3.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a3.operation_mode = "bidir_dual_port";
defparam ram_block3a3.port_a_address_clear = "none";
defparam ram_block3a3.port_a_address_width = 13;
defparam ram_block3a3.port_a_byte_enable_clock = "none";
defparam ram_block3a3.port_a_data_out_clear = "none";
defparam ram_block3a3.port_a_data_out_clock = "none";
defparam ram_block3a3.port_a_data_width = 1;
defparam ram_block3a3.port_a_first_address = 0;
defparam ram_block3a3.port_a_first_bit_number = 3;
defparam ram_block3a3.port_a_last_address = 8191;
defparam ram_block3a3.port_a_logical_ram_depth = 16384;
defparam ram_block3a3.port_a_logical_ram_width = 32;
defparam ram_block3a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_address_clear = "none";
defparam ram_block3a3.port_b_address_clock = "clock1";
defparam ram_block3a3.port_b_address_width = 13;
defparam ram_block3a3.port_b_data_in_clock = "clock1";
defparam ram_block3a3.port_b_data_out_clear = "none";
defparam ram_block3a3.port_b_data_out_clock = "none";
defparam ram_block3a3.port_b_data_width = 1;
defparam ram_block3a3.port_b_first_address = 0;
defparam ram_block3a3.port_b_first_bit_number = 3;
defparam ram_block3a3.port_b_last_address = 8191;
defparam ram_block3a3.port_b_logical_ram_depth = 16384;
defparam ram_block3a3.port_b_logical_ram_width = 32;
defparam ram_block3a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_read_enable_clock = "clock1";
defparam ram_block3a3.port_b_write_enable_clock = "clock1";
defparam ram_block3a3.ram_block_type = "M9K";
defparam ram_block3a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009F20E64C2468E52000000000000000000000000000022346308C62632A08083;
// synopsys translate_on

// Location: M9K_X64_Y42_N0
cycloneive_ram_block ram_block3a36(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a36_PORTADATAOUT_bus),
	.portbdataout(ram_block3a36_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a36.clk0_core_clock_enable = "ena0";
defparam ram_block3a36.clk1_core_clock_enable = "ena1";
defparam ram_block3a36.data_interleave_offset_in_bits = 1;
defparam ram_block3a36.data_interleave_width_in_bits = 1;
defparam ram_block3a36.init_file = "meminit.hex";
defparam ram_block3a36.init_file_layout = "port_a";
defparam ram_block3a36.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a36.operation_mode = "bidir_dual_port";
defparam ram_block3a36.port_a_address_clear = "none";
defparam ram_block3a36.port_a_address_width = 13;
defparam ram_block3a36.port_a_byte_enable_clock = "none";
defparam ram_block3a36.port_a_data_out_clear = "none";
defparam ram_block3a36.port_a_data_out_clock = "none";
defparam ram_block3a36.port_a_data_width = 1;
defparam ram_block3a36.port_a_first_address = 0;
defparam ram_block3a36.port_a_first_bit_number = 4;
defparam ram_block3a36.port_a_last_address = 8191;
defparam ram_block3a36.port_a_logical_ram_depth = 16384;
defparam ram_block3a36.port_a_logical_ram_width = 32;
defparam ram_block3a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_address_clear = "none";
defparam ram_block3a36.port_b_address_clock = "clock1";
defparam ram_block3a36.port_b_address_width = 13;
defparam ram_block3a36.port_b_data_in_clock = "clock1";
defparam ram_block3a36.port_b_data_out_clear = "none";
defparam ram_block3a36.port_b_data_out_clock = "none";
defparam ram_block3a36.port_b_data_width = 1;
defparam ram_block3a36.port_b_first_address = 0;
defparam ram_block3a36.port_b_first_bit_number = 4;
defparam ram_block3a36.port_b_last_address = 8191;
defparam ram_block3a36.port_b_logical_ram_depth = 16384;
defparam ram_block3a36.port_b_logical_ram_width = 32;
defparam ram_block3a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_read_enable_clock = "clock1";
defparam ram_block3a36.port_b_write_enable_clock = "clock1";
defparam ram_block3a36.ram_block_type = "M9K";
defparam ram_block3a36.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y41_N0
cycloneive_ram_block ram_block3a4(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a4_PORTADATAOUT_bus),
	.portbdataout(ram_block3a4_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a4.clk0_core_clock_enable = "ena0";
defparam ram_block3a4.clk1_core_clock_enable = "ena1";
defparam ram_block3a4.data_interleave_offset_in_bits = 1;
defparam ram_block3a4.data_interleave_width_in_bits = 1;
defparam ram_block3a4.init_file = "meminit.hex";
defparam ram_block3a4.init_file_layout = "port_a";
defparam ram_block3a4.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a4.operation_mode = "bidir_dual_port";
defparam ram_block3a4.port_a_address_clear = "none";
defparam ram_block3a4.port_a_address_width = 13;
defparam ram_block3a4.port_a_byte_enable_clock = "none";
defparam ram_block3a4.port_a_data_out_clear = "none";
defparam ram_block3a4.port_a_data_out_clock = "none";
defparam ram_block3a4.port_a_data_width = 1;
defparam ram_block3a4.port_a_first_address = 0;
defparam ram_block3a4.port_a_first_bit_number = 4;
defparam ram_block3a4.port_a_last_address = 8191;
defparam ram_block3a4.port_a_logical_ram_depth = 16384;
defparam ram_block3a4.port_a_logical_ram_width = 32;
defparam ram_block3a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_address_clear = "none";
defparam ram_block3a4.port_b_address_clock = "clock1";
defparam ram_block3a4.port_b_address_width = 13;
defparam ram_block3a4.port_b_data_in_clock = "clock1";
defparam ram_block3a4.port_b_data_out_clear = "none";
defparam ram_block3a4.port_b_data_out_clock = "none";
defparam ram_block3a4.port_b_data_width = 1;
defparam ram_block3a4.port_b_first_address = 0;
defparam ram_block3a4.port_b_first_bit_number = 4;
defparam ram_block3a4.port_b_last_address = 8191;
defparam ram_block3a4.port_b_logical_ram_depth = 16384;
defparam ram_block3a4.port_b_logical_ram_width = 32;
defparam ram_block3a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_read_enable_clock = "clock1";
defparam ram_block3a4.port_b_write_enable_clock = "clock1";
defparam ram_block3a4.ram_block_type = "M9K";
defparam ram_block3a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060B81842D24565BE000000000000000000000000000002242101022202208083;
// synopsys translate_on

// Location: M9K_X51_Y30_N0
cycloneive_ram_block ram_block3a37(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a37_PORTADATAOUT_bus),
	.portbdataout(ram_block3a37_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a37.clk0_core_clock_enable = "ena0";
defparam ram_block3a37.clk1_core_clock_enable = "ena1";
defparam ram_block3a37.data_interleave_offset_in_bits = 1;
defparam ram_block3a37.data_interleave_width_in_bits = 1;
defparam ram_block3a37.init_file = "meminit.hex";
defparam ram_block3a37.init_file_layout = "port_a";
defparam ram_block3a37.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a37.operation_mode = "bidir_dual_port";
defparam ram_block3a37.port_a_address_clear = "none";
defparam ram_block3a37.port_a_address_width = 13;
defparam ram_block3a37.port_a_byte_enable_clock = "none";
defparam ram_block3a37.port_a_data_out_clear = "none";
defparam ram_block3a37.port_a_data_out_clock = "none";
defparam ram_block3a37.port_a_data_width = 1;
defparam ram_block3a37.port_a_first_address = 0;
defparam ram_block3a37.port_a_first_bit_number = 5;
defparam ram_block3a37.port_a_last_address = 8191;
defparam ram_block3a37.port_a_logical_ram_depth = 16384;
defparam ram_block3a37.port_a_logical_ram_width = 32;
defparam ram_block3a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_address_clear = "none";
defparam ram_block3a37.port_b_address_clock = "clock1";
defparam ram_block3a37.port_b_address_width = 13;
defparam ram_block3a37.port_b_data_in_clock = "clock1";
defparam ram_block3a37.port_b_data_out_clear = "none";
defparam ram_block3a37.port_b_data_out_clock = "none";
defparam ram_block3a37.port_b_data_width = 1;
defparam ram_block3a37.port_b_first_address = 0;
defparam ram_block3a37.port_b_first_bit_number = 5;
defparam ram_block3a37.port_b_last_address = 8191;
defparam ram_block3a37.port_b_logical_ram_depth = 16384;
defparam ram_block3a37.port_b_logical_ram_width = 32;
defparam ram_block3a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_read_enable_clock = "clock1";
defparam ram_block3a37.port_b_write_enable_clock = "clock1";
defparam ram_block3a37.ram_block_type = "M9K";
defparam ram_block3a37.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y26_N0
cycloneive_ram_block ram_block3a5(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a5_PORTADATAOUT_bus),
	.portbdataout(ram_block3a5_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a5.clk0_core_clock_enable = "ena0";
defparam ram_block3a5.clk1_core_clock_enable = "ena1";
defparam ram_block3a5.data_interleave_offset_in_bits = 1;
defparam ram_block3a5.data_interleave_width_in_bits = 1;
defparam ram_block3a5.init_file = "meminit.hex";
defparam ram_block3a5.init_file_layout = "port_a";
defparam ram_block3a5.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a5.operation_mode = "bidir_dual_port";
defparam ram_block3a5.port_a_address_clear = "none";
defparam ram_block3a5.port_a_address_width = 13;
defparam ram_block3a5.port_a_byte_enable_clock = "none";
defparam ram_block3a5.port_a_data_out_clear = "none";
defparam ram_block3a5.port_a_data_out_clock = "none";
defparam ram_block3a5.port_a_data_width = 1;
defparam ram_block3a5.port_a_first_address = 0;
defparam ram_block3a5.port_a_first_bit_number = 5;
defparam ram_block3a5.port_a_last_address = 8191;
defparam ram_block3a5.port_a_logical_ram_depth = 16384;
defparam ram_block3a5.port_a_logical_ram_width = 32;
defparam ram_block3a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_address_clear = "none";
defparam ram_block3a5.port_b_address_clock = "clock1";
defparam ram_block3a5.port_b_address_width = 13;
defparam ram_block3a5.port_b_data_in_clock = "clock1";
defparam ram_block3a5.port_b_data_out_clear = "none";
defparam ram_block3a5.port_b_data_out_clock = "none";
defparam ram_block3a5.port_b_data_width = 1;
defparam ram_block3a5.port_b_first_address = 0;
defparam ram_block3a5.port_b_first_bit_number = 5;
defparam ram_block3a5.port_b_last_address = 8191;
defparam ram_block3a5.port_b_logical_ram_depth = 16384;
defparam ram_block3a5.port_b_logical_ram_width = 32;
defparam ram_block3a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_read_enable_clock = "clock1";
defparam ram_block3a5.port_b_write_enable_clock = "clock1";
defparam ram_block3a5.ram_block_type = "M9K";
defparam ram_block3a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000056414512D6B00448000000000000000000000000000002246308006652AF7263;
// synopsys translate_on

// Location: M9K_X64_Y27_N0
cycloneive_ram_block ram_block3a38(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a38_PORTADATAOUT_bus),
	.portbdataout(ram_block3a38_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a38.clk0_core_clock_enable = "ena0";
defparam ram_block3a38.clk1_core_clock_enable = "ena1";
defparam ram_block3a38.data_interleave_offset_in_bits = 1;
defparam ram_block3a38.data_interleave_width_in_bits = 1;
defparam ram_block3a38.init_file = "meminit.hex";
defparam ram_block3a38.init_file_layout = "port_a";
defparam ram_block3a38.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a38.operation_mode = "bidir_dual_port";
defparam ram_block3a38.port_a_address_clear = "none";
defparam ram_block3a38.port_a_address_width = 13;
defparam ram_block3a38.port_a_byte_enable_clock = "none";
defparam ram_block3a38.port_a_data_out_clear = "none";
defparam ram_block3a38.port_a_data_out_clock = "none";
defparam ram_block3a38.port_a_data_width = 1;
defparam ram_block3a38.port_a_first_address = 0;
defparam ram_block3a38.port_a_first_bit_number = 6;
defparam ram_block3a38.port_a_last_address = 8191;
defparam ram_block3a38.port_a_logical_ram_depth = 16384;
defparam ram_block3a38.port_a_logical_ram_width = 32;
defparam ram_block3a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_address_clear = "none";
defparam ram_block3a38.port_b_address_clock = "clock1";
defparam ram_block3a38.port_b_address_width = 13;
defparam ram_block3a38.port_b_data_in_clock = "clock1";
defparam ram_block3a38.port_b_data_out_clear = "none";
defparam ram_block3a38.port_b_data_out_clock = "none";
defparam ram_block3a38.port_b_data_width = 1;
defparam ram_block3a38.port_b_first_address = 0;
defparam ram_block3a38.port_b_first_bit_number = 6;
defparam ram_block3a38.port_b_last_address = 8191;
defparam ram_block3a38.port_b_logical_ram_depth = 16384;
defparam ram_block3a38.port_b_logical_ram_width = 32;
defparam ram_block3a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_read_enable_clock = "clock1";
defparam ram_block3a38.port_b_write_enable_clock = "clock1";
defparam ram_block3a38.ram_block_type = "M9K";
defparam ram_block3a38.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y30_N0
cycloneive_ram_block ram_block3a6(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a6_PORTADATAOUT_bus),
	.portbdataout(ram_block3a6_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a6.clk0_core_clock_enable = "ena0";
defparam ram_block3a6.clk1_core_clock_enable = "ena1";
defparam ram_block3a6.data_interleave_offset_in_bits = 1;
defparam ram_block3a6.data_interleave_width_in_bits = 1;
defparam ram_block3a6.init_file = "meminit.hex";
defparam ram_block3a6.init_file_layout = "port_a";
defparam ram_block3a6.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a6.operation_mode = "bidir_dual_port";
defparam ram_block3a6.port_a_address_clear = "none";
defparam ram_block3a6.port_a_address_width = 13;
defparam ram_block3a6.port_a_byte_enable_clock = "none";
defparam ram_block3a6.port_a_data_out_clear = "none";
defparam ram_block3a6.port_a_data_out_clock = "none";
defparam ram_block3a6.port_a_data_width = 1;
defparam ram_block3a6.port_a_first_address = 0;
defparam ram_block3a6.port_a_first_bit_number = 6;
defparam ram_block3a6.port_a_last_address = 8191;
defparam ram_block3a6.port_a_logical_ram_depth = 16384;
defparam ram_block3a6.port_a_logical_ram_width = 32;
defparam ram_block3a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_address_clear = "none";
defparam ram_block3a6.port_b_address_clock = "clock1";
defparam ram_block3a6.port_b_address_width = 13;
defparam ram_block3a6.port_b_data_in_clock = "clock1";
defparam ram_block3a6.port_b_data_out_clear = "none";
defparam ram_block3a6.port_b_data_out_clock = "none";
defparam ram_block3a6.port_b_data_width = 1;
defparam ram_block3a6.port_b_first_address = 0;
defparam ram_block3a6.port_b_first_bit_number = 6;
defparam ram_block3a6.port_b_last_address = 8191;
defparam ram_block3a6.port_b_logical_ram_depth = 16384;
defparam ram_block3a6.port_b_logical_ram_width = 32;
defparam ram_block3a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_read_enable_clock = "clock1";
defparam ram_block3a6.port_b_write_enable_clock = "clock1";
defparam ram_block3a6.ram_block_type = "M9K";
defparam ram_block3a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001003088D801A0F827000000000000000000000000000012042100402202200113;
// synopsys translate_on

// Location: M9K_X51_Y42_N0
cycloneive_ram_block ram_block3a39(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a39_PORTADATAOUT_bus),
	.portbdataout(ram_block3a39_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a39.clk0_core_clock_enable = "ena0";
defparam ram_block3a39.clk1_core_clock_enable = "ena1";
defparam ram_block3a39.data_interleave_offset_in_bits = 1;
defparam ram_block3a39.data_interleave_width_in_bits = 1;
defparam ram_block3a39.init_file = "meminit.hex";
defparam ram_block3a39.init_file_layout = "port_a";
defparam ram_block3a39.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a39.operation_mode = "bidir_dual_port";
defparam ram_block3a39.port_a_address_clear = "none";
defparam ram_block3a39.port_a_address_width = 13;
defparam ram_block3a39.port_a_byte_enable_clock = "none";
defparam ram_block3a39.port_a_data_out_clear = "none";
defparam ram_block3a39.port_a_data_out_clock = "none";
defparam ram_block3a39.port_a_data_width = 1;
defparam ram_block3a39.port_a_first_address = 0;
defparam ram_block3a39.port_a_first_bit_number = 7;
defparam ram_block3a39.port_a_last_address = 8191;
defparam ram_block3a39.port_a_logical_ram_depth = 16384;
defparam ram_block3a39.port_a_logical_ram_width = 32;
defparam ram_block3a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_address_clear = "none";
defparam ram_block3a39.port_b_address_clock = "clock1";
defparam ram_block3a39.port_b_address_width = 13;
defparam ram_block3a39.port_b_data_in_clock = "clock1";
defparam ram_block3a39.port_b_data_out_clear = "none";
defparam ram_block3a39.port_b_data_out_clock = "none";
defparam ram_block3a39.port_b_data_width = 1;
defparam ram_block3a39.port_b_first_address = 0;
defparam ram_block3a39.port_b_first_bit_number = 7;
defparam ram_block3a39.port_b_last_address = 8191;
defparam ram_block3a39.port_b_logical_ram_depth = 16384;
defparam ram_block3a39.port_b_logical_ram_width = 32;
defparam ram_block3a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_read_enable_clock = "clock1";
defparam ram_block3a39.port_b_write_enable_clock = "clock1";
defparam ram_block3a39.ram_block_type = "M9K";
defparam ram_block3a39.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y40_N0
cycloneive_ram_block ram_block3a7(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a7_PORTADATAOUT_bus),
	.portbdataout(ram_block3a7_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a7.clk0_core_clock_enable = "ena0";
defparam ram_block3a7.clk1_core_clock_enable = "ena1";
defparam ram_block3a7.data_interleave_offset_in_bits = 1;
defparam ram_block3a7.data_interleave_width_in_bits = 1;
defparam ram_block3a7.init_file = "meminit.hex";
defparam ram_block3a7.init_file_layout = "port_a";
defparam ram_block3a7.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a7.operation_mode = "bidir_dual_port";
defparam ram_block3a7.port_a_address_clear = "none";
defparam ram_block3a7.port_a_address_width = 13;
defparam ram_block3a7.port_a_byte_enable_clock = "none";
defparam ram_block3a7.port_a_data_out_clear = "none";
defparam ram_block3a7.port_a_data_out_clock = "none";
defparam ram_block3a7.port_a_data_width = 1;
defparam ram_block3a7.port_a_first_address = 0;
defparam ram_block3a7.port_a_first_bit_number = 7;
defparam ram_block3a7.port_a_last_address = 8191;
defparam ram_block3a7.port_a_logical_ram_depth = 16384;
defparam ram_block3a7.port_a_logical_ram_width = 32;
defparam ram_block3a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_address_clear = "none";
defparam ram_block3a7.port_b_address_clock = "clock1";
defparam ram_block3a7.port_b_address_width = 13;
defparam ram_block3a7.port_b_data_in_clock = "clock1";
defparam ram_block3a7.port_b_data_out_clear = "none";
defparam ram_block3a7.port_b_data_out_clock = "none";
defparam ram_block3a7.port_b_data_width = 1;
defparam ram_block3a7.port_b_first_address = 0;
defparam ram_block3a7.port_b_first_bit_number = 7;
defparam ram_block3a7.port_b_last_address = 8191;
defparam ram_block3a7.port_b_logical_ram_depth = 16384;
defparam ram_block3a7.port_b_logical_ram_width = 32;
defparam ram_block3a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_read_enable_clock = "clock1";
defparam ram_block3a7.port_b_write_enable_clock = "clock1";
defparam ram_block3a7.ram_block_type = "M9K";
defparam ram_block3a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220A200403;
// synopsys translate_on

// Location: M9K_X51_Y34_N0
cycloneive_ram_block ram_block3a40(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a40_PORTADATAOUT_bus),
	.portbdataout(ram_block3a40_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a40.clk0_core_clock_enable = "ena0";
defparam ram_block3a40.clk1_core_clock_enable = "ena1";
defparam ram_block3a40.data_interleave_offset_in_bits = 1;
defparam ram_block3a40.data_interleave_width_in_bits = 1;
defparam ram_block3a40.init_file = "meminit.hex";
defparam ram_block3a40.init_file_layout = "port_a";
defparam ram_block3a40.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a40.operation_mode = "bidir_dual_port";
defparam ram_block3a40.port_a_address_clear = "none";
defparam ram_block3a40.port_a_address_width = 13;
defparam ram_block3a40.port_a_byte_enable_clock = "none";
defparam ram_block3a40.port_a_data_out_clear = "none";
defparam ram_block3a40.port_a_data_out_clock = "none";
defparam ram_block3a40.port_a_data_width = 1;
defparam ram_block3a40.port_a_first_address = 0;
defparam ram_block3a40.port_a_first_bit_number = 8;
defparam ram_block3a40.port_a_last_address = 8191;
defparam ram_block3a40.port_a_logical_ram_depth = 16384;
defparam ram_block3a40.port_a_logical_ram_width = 32;
defparam ram_block3a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_address_clear = "none";
defparam ram_block3a40.port_b_address_clock = "clock1";
defparam ram_block3a40.port_b_address_width = 13;
defparam ram_block3a40.port_b_data_in_clock = "clock1";
defparam ram_block3a40.port_b_data_out_clear = "none";
defparam ram_block3a40.port_b_data_out_clock = "none";
defparam ram_block3a40.port_b_data_width = 1;
defparam ram_block3a40.port_b_first_address = 0;
defparam ram_block3a40.port_b_first_bit_number = 8;
defparam ram_block3a40.port_b_last_address = 8191;
defparam ram_block3a40.port_b_logical_ram_depth = 16384;
defparam ram_block3a40.port_b_logical_ram_width = 32;
defparam ram_block3a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_read_enable_clock = "clock1";
defparam ram_block3a40.port_b_write_enable_clock = "clock1";
defparam ram_block3a40.ram_block_type = "M9K";
defparam ram_block3a40.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y34_N0
cycloneive_ram_block ram_block3a8(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a8_PORTADATAOUT_bus),
	.portbdataout(ram_block3a8_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a8.clk0_core_clock_enable = "ena0";
defparam ram_block3a8.clk1_core_clock_enable = "ena1";
defparam ram_block3a8.data_interleave_offset_in_bits = 1;
defparam ram_block3a8.data_interleave_width_in_bits = 1;
defparam ram_block3a8.init_file = "meminit.hex";
defparam ram_block3a8.init_file_layout = "port_a";
defparam ram_block3a8.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a8.operation_mode = "bidir_dual_port";
defparam ram_block3a8.port_a_address_clear = "none";
defparam ram_block3a8.port_a_address_width = 13;
defparam ram_block3a8.port_a_byte_enable_clock = "none";
defparam ram_block3a8.port_a_data_out_clear = "none";
defparam ram_block3a8.port_a_data_out_clock = "none";
defparam ram_block3a8.port_a_data_width = 1;
defparam ram_block3a8.port_a_first_address = 0;
defparam ram_block3a8.port_a_first_bit_number = 8;
defparam ram_block3a8.port_a_last_address = 8191;
defparam ram_block3a8.port_a_logical_ram_depth = 16384;
defparam ram_block3a8.port_a_logical_ram_width = 32;
defparam ram_block3a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_address_clear = "none";
defparam ram_block3a8.port_b_address_clock = "clock1";
defparam ram_block3a8.port_b_address_width = 13;
defparam ram_block3a8.port_b_data_in_clock = "clock1";
defparam ram_block3a8.port_b_data_out_clear = "none";
defparam ram_block3a8.port_b_data_out_clock = "none";
defparam ram_block3a8.port_b_data_width = 1;
defparam ram_block3a8.port_b_first_address = 0;
defparam ram_block3a8.port_b_first_bit_number = 8;
defparam ram_block3a8.port_b_last_address = 8191;
defparam ram_block3a8.port_b_logical_ram_depth = 16384;
defparam ram_block3a8.port_b_logical_ram_width = 32;
defparam ram_block3a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_read_enable_clock = "clock1";
defparam ram_block3a8.port_b_write_enable_clock = "clock1";
defparam ram_block3a8.ram_block_type = "M9K";
defparam ram_block3a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220230080F;
// synopsys translate_on

// Location: M9K_X78_Y38_N0
cycloneive_ram_block ram_block3a41(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a41_PORTADATAOUT_bus),
	.portbdataout(ram_block3a41_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a41.clk0_core_clock_enable = "ena0";
defparam ram_block3a41.clk1_core_clock_enable = "ena1";
defparam ram_block3a41.data_interleave_offset_in_bits = 1;
defparam ram_block3a41.data_interleave_width_in_bits = 1;
defparam ram_block3a41.init_file = "meminit.hex";
defparam ram_block3a41.init_file_layout = "port_a";
defparam ram_block3a41.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a41.operation_mode = "bidir_dual_port";
defparam ram_block3a41.port_a_address_clear = "none";
defparam ram_block3a41.port_a_address_width = 13;
defparam ram_block3a41.port_a_byte_enable_clock = "none";
defparam ram_block3a41.port_a_data_out_clear = "none";
defparam ram_block3a41.port_a_data_out_clock = "none";
defparam ram_block3a41.port_a_data_width = 1;
defparam ram_block3a41.port_a_first_address = 0;
defparam ram_block3a41.port_a_first_bit_number = 9;
defparam ram_block3a41.port_a_last_address = 8191;
defparam ram_block3a41.port_a_logical_ram_depth = 16384;
defparam ram_block3a41.port_a_logical_ram_width = 32;
defparam ram_block3a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_address_clear = "none";
defparam ram_block3a41.port_b_address_clock = "clock1";
defparam ram_block3a41.port_b_address_width = 13;
defparam ram_block3a41.port_b_data_in_clock = "clock1";
defparam ram_block3a41.port_b_data_out_clear = "none";
defparam ram_block3a41.port_b_data_out_clock = "none";
defparam ram_block3a41.port_b_data_width = 1;
defparam ram_block3a41.port_b_first_address = 0;
defparam ram_block3a41.port_b_first_bit_number = 9;
defparam ram_block3a41.port_b_last_address = 8191;
defparam ram_block3a41.port_b_logical_ram_depth = 16384;
defparam ram_block3a41.port_b_logical_ram_width = 32;
defparam ram_block3a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_read_enable_clock = "clock1";
defparam ram_block3a41.port_b_write_enable_clock = "clock1";
defparam ram_block3a41.ram_block_type = "M9K";
defparam ram_block3a41.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y40_N0
cycloneive_ram_block ram_block3a9(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a9_PORTADATAOUT_bus),
	.portbdataout(ram_block3a9_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a9.clk0_core_clock_enable = "ena0";
defparam ram_block3a9.clk1_core_clock_enable = "ena1";
defparam ram_block3a9.data_interleave_offset_in_bits = 1;
defparam ram_block3a9.data_interleave_width_in_bits = 1;
defparam ram_block3a9.init_file = "meminit.hex";
defparam ram_block3a9.init_file_layout = "port_a";
defparam ram_block3a9.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a9.operation_mode = "bidir_dual_port";
defparam ram_block3a9.port_a_address_clear = "none";
defparam ram_block3a9.port_a_address_width = 13;
defparam ram_block3a9.port_a_byte_enable_clock = "none";
defparam ram_block3a9.port_a_data_out_clear = "none";
defparam ram_block3a9.port_a_data_out_clock = "none";
defparam ram_block3a9.port_a_data_width = 1;
defparam ram_block3a9.port_a_first_address = 0;
defparam ram_block3a9.port_a_first_bit_number = 9;
defparam ram_block3a9.port_a_last_address = 8191;
defparam ram_block3a9.port_a_logical_ram_depth = 16384;
defparam ram_block3a9.port_a_logical_ram_width = 32;
defparam ram_block3a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_address_clear = "none";
defparam ram_block3a9.port_b_address_clock = "clock1";
defparam ram_block3a9.port_b_address_width = 13;
defparam ram_block3a9.port_b_data_in_clock = "clock1";
defparam ram_block3a9.port_b_data_out_clear = "none";
defparam ram_block3a9.port_b_data_out_clock = "none";
defparam ram_block3a9.port_b_data_width = 1;
defparam ram_block3a9.port_b_first_address = 0;
defparam ram_block3a9.port_b_first_bit_number = 9;
defparam ram_block3a9.port_b_last_address = 8191;
defparam ram_block3a9.port_b_logical_ram_depth = 16384;
defparam ram_block3a9.port_b_logical_ram_width = 32;
defparam ram_block3a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_read_enable_clock = "clock1";
defparam ram_block3a9.port_b_write_enable_clock = "clock1";
defparam ram_block3a9.ram_block_type = "M9K";
defparam ram_block3a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220220080F;
// synopsys translate_on

// Location: M9K_X51_Y38_N0
cycloneive_ram_block ram_block3a42(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a42_PORTADATAOUT_bus),
	.portbdataout(ram_block3a42_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a42.clk0_core_clock_enable = "ena0";
defparam ram_block3a42.clk1_core_clock_enable = "ena1";
defparam ram_block3a42.data_interleave_offset_in_bits = 1;
defparam ram_block3a42.data_interleave_width_in_bits = 1;
defparam ram_block3a42.init_file = "meminit.hex";
defparam ram_block3a42.init_file_layout = "port_a";
defparam ram_block3a42.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a42.operation_mode = "bidir_dual_port";
defparam ram_block3a42.port_a_address_clear = "none";
defparam ram_block3a42.port_a_address_width = 13;
defparam ram_block3a42.port_a_byte_enable_clock = "none";
defparam ram_block3a42.port_a_data_out_clear = "none";
defparam ram_block3a42.port_a_data_out_clock = "none";
defparam ram_block3a42.port_a_data_width = 1;
defparam ram_block3a42.port_a_first_address = 0;
defparam ram_block3a42.port_a_first_bit_number = 10;
defparam ram_block3a42.port_a_last_address = 8191;
defparam ram_block3a42.port_a_logical_ram_depth = 16384;
defparam ram_block3a42.port_a_logical_ram_width = 32;
defparam ram_block3a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_address_clear = "none";
defparam ram_block3a42.port_b_address_clock = "clock1";
defparam ram_block3a42.port_b_address_width = 13;
defparam ram_block3a42.port_b_data_in_clock = "clock1";
defparam ram_block3a42.port_b_data_out_clear = "none";
defparam ram_block3a42.port_b_data_out_clock = "none";
defparam ram_block3a42.port_b_data_width = 1;
defparam ram_block3a42.port_b_first_address = 0;
defparam ram_block3a42.port_b_first_bit_number = 10;
defparam ram_block3a42.port_b_last_address = 8191;
defparam ram_block3a42.port_b_logical_ram_depth = 16384;
defparam ram_block3a42.port_b_logical_ram_width = 32;
defparam ram_block3a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_read_enable_clock = "clock1";
defparam ram_block3a42.port_b_write_enable_clock = "clock1";
defparam ram_block3a42.ram_block_type = "M9K";
defparam ram_block3a42.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y38_N0
cycloneive_ram_block ram_block3a10(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a10_PORTADATAOUT_bus),
	.portbdataout(ram_block3a10_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a10.clk0_core_clock_enable = "ena0";
defparam ram_block3a10.clk1_core_clock_enable = "ena1";
defparam ram_block3a10.data_interleave_offset_in_bits = 1;
defparam ram_block3a10.data_interleave_width_in_bits = 1;
defparam ram_block3a10.init_file = "meminit.hex";
defparam ram_block3a10.init_file_layout = "port_a";
defparam ram_block3a10.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a10.operation_mode = "bidir_dual_port";
defparam ram_block3a10.port_a_address_clear = "none";
defparam ram_block3a10.port_a_address_width = 13;
defparam ram_block3a10.port_a_byte_enable_clock = "none";
defparam ram_block3a10.port_a_data_out_clear = "none";
defparam ram_block3a10.port_a_data_out_clock = "none";
defparam ram_block3a10.port_a_data_width = 1;
defparam ram_block3a10.port_a_first_address = 0;
defparam ram_block3a10.port_a_first_bit_number = 10;
defparam ram_block3a10.port_a_last_address = 8191;
defparam ram_block3a10.port_a_logical_ram_depth = 16384;
defparam ram_block3a10.port_a_logical_ram_width = 32;
defparam ram_block3a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_address_clear = "none";
defparam ram_block3a10.port_b_address_clock = "clock1";
defparam ram_block3a10.port_b_address_width = 13;
defparam ram_block3a10.port_b_data_in_clock = "clock1";
defparam ram_block3a10.port_b_data_out_clear = "none";
defparam ram_block3a10.port_b_data_out_clock = "none";
defparam ram_block3a10.port_b_data_width = 1;
defparam ram_block3a10.port_b_first_address = 0;
defparam ram_block3a10.port_b_first_bit_number = 10;
defparam ram_block3a10.port_b_last_address = 8191;
defparam ram_block3a10.port_b_logical_ram_depth = 16384;
defparam ram_block3a10.port_b_logical_ram_width = 32;
defparam ram_block3a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_read_enable_clock = "clock1";
defparam ram_block3a10.port_b_write_enable_clock = "clock1";
defparam ram_block3a10.ram_block_type = "M9K";
defparam ram_block3a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002042100002202300003;
// synopsys translate_on

// Location: M9K_X51_Y32_N0
cycloneive_ram_block ram_block3a43(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a43_PORTADATAOUT_bus),
	.portbdataout(ram_block3a43_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a43.clk0_core_clock_enable = "ena0";
defparam ram_block3a43.clk1_core_clock_enable = "ena1";
defparam ram_block3a43.data_interleave_offset_in_bits = 1;
defparam ram_block3a43.data_interleave_width_in_bits = 1;
defparam ram_block3a43.init_file = "meminit.hex";
defparam ram_block3a43.init_file_layout = "port_a";
defparam ram_block3a43.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a43.operation_mode = "bidir_dual_port";
defparam ram_block3a43.port_a_address_clear = "none";
defparam ram_block3a43.port_a_address_width = 13;
defparam ram_block3a43.port_a_byte_enable_clock = "none";
defparam ram_block3a43.port_a_data_out_clear = "none";
defparam ram_block3a43.port_a_data_out_clock = "none";
defparam ram_block3a43.port_a_data_width = 1;
defparam ram_block3a43.port_a_first_address = 0;
defparam ram_block3a43.port_a_first_bit_number = 11;
defparam ram_block3a43.port_a_last_address = 8191;
defparam ram_block3a43.port_a_logical_ram_depth = 16384;
defparam ram_block3a43.port_a_logical_ram_width = 32;
defparam ram_block3a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_address_clear = "none";
defparam ram_block3a43.port_b_address_clock = "clock1";
defparam ram_block3a43.port_b_address_width = 13;
defparam ram_block3a43.port_b_data_in_clock = "clock1";
defparam ram_block3a43.port_b_data_out_clear = "none";
defparam ram_block3a43.port_b_data_out_clock = "none";
defparam ram_block3a43.port_b_data_width = 1;
defparam ram_block3a43.port_b_first_address = 0;
defparam ram_block3a43.port_b_first_bit_number = 11;
defparam ram_block3a43.port_b_last_address = 8191;
defparam ram_block3a43.port_b_logical_ram_depth = 16384;
defparam ram_block3a43.port_b_logical_ram_width = 32;
defparam ram_block3a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_read_enable_clock = "clock1";
defparam ram_block3a43.port_b_write_enable_clock = "clock1";
defparam ram_block3a43.ram_block_type = "M9K";
defparam ram_block3a43.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y31_N0
cycloneive_ram_block ram_block3a11(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a11_PORTADATAOUT_bus),
	.portbdataout(ram_block3a11_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a11.clk0_core_clock_enable = "ena0";
defparam ram_block3a11.clk1_core_clock_enable = "ena1";
defparam ram_block3a11.data_interleave_offset_in_bits = 1;
defparam ram_block3a11.data_interleave_width_in_bits = 1;
defparam ram_block3a11.init_file = "meminit.hex";
defparam ram_block3a11.init_file_layout = "port_a";
defparam ram_block3a11.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a11.operation_mode = "bidir_dual_port";
defparam ram_block3a11.port_a_address_clear = "none";
defparam ram_block3a11.port_a_address_width = 13;
defparam ram_block3a11.port_a_byte_enable_clock = "none";
defparam ram_block3a11.port_a_data_out_clear = "none";
defparam ram_block3a11.port_a_data_out_clock = "none";
defparam ram_block3a11.port_a_data_width = 1;
defparam ram_block3a11.port_a_first_address = 0;
defparam ram_block3a11.port_a_first_bit_number = 11;
defparam ram_block3a11.port_a_last_address = 8191;
defparam ram_block3a11.port_a_logical_ram_depth = 16384;
defparam ram_block3a11.port_a_logical_ram_width = 32;
defparam ram_block3a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_address_clear = "none";
defparam ram_block3a11.port_b_address_clock = "clock1";
defparam ram_block3a11.port_b_address_width = 13;
defparam ram_block3a11.port_b_data_in_clock = "clock1";
defparam ram_block3a11.port_b_data_out_clear = "none";
defparam ram_block3a11.port_b_data_out_clock = "none";
defparam ram_block3a11.port_b_data_width = 1;
defparam ram_block3a11.port_b_first_address = 0;
defparam ram_block3a11.port_b_first_bit_number = 11;
defparam ram_block3a11.port_b_last_address = 8191;
defparam ram_block3a11.port_b_logical_ram_depth = 16384;
defparam ram_block3a11.port_b_logical_ram_width = 32;
defparam ram_block3a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_read_enable_clock = "clock1";
defparam ram_block3a11.port_b_write_enable_clock = "clock1";
defparam ram_block3a11.ram_block_type = "M9K";
defparam ram_block3a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210800265A2A2233;
// synopsys translate_on

// Location: M9K_X64_Y35_N0
cycloneive_ram_block ram_block3a44(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a44_PORTADATAOUT_bus),
	.portbdataout(ram_block3a44_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a44.clk0_core_clock_enable = "ena0";
defparam ram_block3a44.clk1_core_clock_enable = "ena1";
defparam ram_block3a44.data_interleave_offset_in_bits = 1;
defparam ram_block3a44.data_interleave_width_in_bits = 1;
defparam ram_block3a44.init_file = "meminit.hex";
defparam ram_block3a44.init_file_layout = "port_a";
defparam ram_block3a44.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a44.operation_mode = "bidir_dual_port";
defparam ram_block3a44.port_a_address_clear = "none";
defparam ram_block3a44.port_a_address_width = 13;
defparam ram_block3a44.port_a_byte_enable_clock = "none";
defparam ram_block3a44.port_a_data_out_clear = "none";
defparam ram_block3a44.port_a_data_out_clock = "none";
defparam ram_block3a44.port_a_data_width = 1;
defparam ram_block3a44.port_a_first_address = 0;
defparam ram_block3a44.port_a_first_bit_number = 12;
defparam ram_block3a44.port_a_last_address = 8191;
defparam ram_block3a44.port_a_logical_ram_depth = 16384;
defparam ram_block3a44.port_a_logical_ram_width = 32;
defparam ram_block3a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_address_clear = "none";
defparam ram_block3a44.port_b_address_clock = "clock1";
defparam ram_block3a44.port_b_address_width = 13;
defparam ram_block3a44.port_b_data_in_clock = "clock1";
defparam ram_block3a44.port_b_data_out_clear = "none";
defparam ram_block3a44.port_b_data_out_clock = "none";
defparam ram_block3a44.port_b_data_width = 1;
defparam ram_block3a44.port_b_first_address = 0;
defparam ram_block3a44.port_b_first_bit_number = 12;
defparam ram_block3a44.port_b_last_address = 8191;
defparam ram_block3a44.port_b_logical_ram_depth = 16384;
defparam ram_block3a44.port_b_logical_ram_width = 32;
defparam ram_block3a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_read_enable_clock = "clock1";
defparam ram_block3a44.port_b_write_enable_clock = "clock1";
defparam ram_block3a44.ram_block_type = "M9K";
defparam ram_block3a44.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y32_N0
cycloneive_ram_block ram_block3a12(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a12_PORTADATAOUT_bus),
	.portbdataout(ram_block3a12_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a12.clk0_core_clock_enable = "ena0";
defparam ram_block3a12.clk1_core_clock_enable = "ena1";
defparam ram_block3a12.data_interleave_offset_in_bits = 1;
defparam ram_block3a12.data_interleave_width_in_bits = 1;
defparam ram_block3a12.init_file = "meminit.hex";
defparam ram_block3a12.init_file_layout = "port_a";
defparam ram_block3a12.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a12.operation_mode = "bidir_dual_port";
defparam ram_block3a12.port_a_address_clear = "none";
defparam ram_block3a12.port_a_address_width = 13;
defparam ram_block3a12.port_a_byte_enable_clock = "none";
defparam ram_block3a12.port_a_data_out_clear = "none";
defparam ram_block3a12.port_a_data_out_clock = "none";
defparam ram_block3a12.port_a_data_width = 1;
defparam ram_block3a12.port_a_first_address = 0;
defparam ram_block3a12.port_a_first_bit_number = 12;
defparam ram_block3a12.port_a_last_address = 8191;
defparam ram_block3a12.port_a_logical_ram_depth = 16384;
defparam ram_block3a12.port_a_logical_ram_width = 32;
defparam ram_block3a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_address_clear = "none";
defparam ram_block3a12.port_b_address_clock = "clock1";
defparam ram_block3a12.port_b_address_width = 13;
defparam ram_block3a12.port_b_data_in_clock = "clock1";
defparam ram_block3a12.port_b_data_out_clear = "none";
defparam ram_block3a12.port_b_data_out_clock = "none";
defparam ram_block3a12.port_b_data_width = 1;
defparam ram_block3a12.port_b_first_address = 0;
defparam ram_block3a12.port_b_first_bit_number = 12;
defparam ram_block3a12.port_b_last_address = 8191;
defparam ram_block3a12.port_b_logical_ram_depth = 16384;
defparam ram_block3a12.port_b_logical_ram_width = 32;
defparam ram_block3a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_read_enable_clock = "clock1";
defparam ram_block3a12.port_b_write_enable_clock = "clock1";
defparam ram_block3a12.ram_block_type = "M9K";
defparam ram_block3a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020421000022022C2043;
// synopsys translate_on

// Location: M9K_X37_Y40_N0
cycloneive_ram_block ram_block3a45(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a45_PORTADATAOUT_bus),
	.portbdataout(ram_block3a45_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a45.clk0_core_clock_enable = "ena0";
defparam ram_block3a45.clk1_core_clock_enable = "ena1";
defparam ram_block3a45.data_interleave_offset_in_bits = 1;
defparam ram_block3a45.data_interleave_width_in_bits = 1;
defparam ram_block3a45.init_file = "meminit.hex";
defparam ram_block3a45.init_file_layout = "port_a";
defparam ram_block3a45.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a45.operation_mode = "bidir_dual_port";
defparam ram_block3a45.port_a_address_clear = "none";
defparam ram_block3a45.port_a_address_width = 13;
defparam ram_block3a45.port_a_byte_enable_clock = "none";
defparam ram_block3a45.port_a_data_out_clear = "none";
defparam ram_block3a45.port_a_data_out_clock = "none";
defparam ram_block3a45.port_a_data_width = 1;
defparam ram_block3a45.port_a_first_address = 0;
defparam ram_block3a45.port_a_first_bit_number = 13;
defparam ram_block3a45.port_a_last_address = 8191;
defparam ram_block3a45.port_a_logical_ram_depth = 16384;
defparam ram_block3a45.port_a_logical_ram_width = 32;
defparam ram_block3a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_address_clear = "none";
defparam ram_block3a45.port_b_address_clock = "clock1";
defparam ram_block3a45.port_b_address_width = 13;
defparam ram_block3a45.port_b_data_in_clock = "clock1";
defparam ram_block3a45.port_b_data_out_clear = "none";
defparam ram_block3a45.port_b_data_out_clock = "none";
defparam ram_block3a45.port_b_data_width = 1;
defparam ram_block3a45.port_b_first_address = 0;
defparam ram_block3a45.port_b_first_bit_number = 13;
defparam ram_block3a45.port_b_last_address = 8191;
defparam ram_block3a45.port_b_logical_ram_depth = 16384;
defparam ram_block3a45.port_b_logical_ram_width = 32;
defparam ram_block3a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_read_enable_clock = "clock1";
defparam ram_block3a45.port_b_write_enable_clock = "clock1";
defparam ram_block3a45.ram_block_type = "M9K";
defparam ram_block3a45.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y41_N0
cycloneive_ram_block ram_block3a13(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a13_PORTADATAOUT_bus),
	.portbdataout(ram_block3a13_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a13.clk0_core_clock_enable = "ena0";
defparam ram_block3a13.clk1_core_clock_enable = "ena1";
defparam ram_block3a13.data_interleave_offset_in_bits = 1;
defparam ram_block3a13.data_interleave_width_in_bits = 1;
defparam ram_block3a13.init_file = "meminit.hex";
defparam ram_block3a13.init_file_layout = "port_a";
defparam ram_block3a13.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a13.operation_mode = "bidir_dual_port";
defparam ram_block3a13.port_a_address_clear = "none";
defparam ram_block3a13.port_a_address_width = 13;
defparam ram_block3a13.port_a_byte_enable_clock = "none";
defparam ram_block3a13.port_a_data_out_clear = "none";
defparam ram_block3a13.port_a_data_out_clock = "none";
defparam ram_block3a13.port_a_data_width = 1;
defparam ram_block3a13.port_a_first_address = 0;
defparam ram_block3a13.port_a_first_bit_number = 13;
defparam ram_block3a13.port_a_last_address = 8191;
defparam ram_block3a13.port_a_logical_ram_depth = 16384;
defparam ram_block3a13.port_a_logical_ram_width = 32;
defparam ram_block3a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_address_clear = "none";
defparam ram_block3a13.port_b_address_clock = "clock1";
defparam ram_block3a13.port_b_address_width = 13;
defparam ram_block3a13.port_b_data_in_clock = "clock1";
defparam ram_block3a13.port_b_data_out_clear = "none";
defparam ram_block3a13.port_b_data_out_clock = "none";
defparam ram_block3a13.port_b_data_width = 1;
defparam ram_block3a13.port_b_first_address = 0;
defparam ram_block3a13.port_b_first_bit_number = 13;
defparam ram_block3a13.port_b_last_address = 8191;
defparam ram_block3a13.port_b_logical_ram_depth = 16384;
defparam ram_block3a13.port_b_logical_ram_width = 32;
defparam ram_block3a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_read_enable_clock = "clock1";
defparam ram_block3a13.port_b_write_enable_clock = "clock1";
defparam ram_block3a13.ram_block_type = "M9K";
defparam ram_block3a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020421000022022F5213;
// synopsys translate_on

// Location: M9K_X37_Y31_N0
cycloneive_ram_block ram_block3a46(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a46_PORTADATAOUT_bus),
	.portbdataout(ram_block3a46_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a46.clk0_core_clock_enable = "ena0";
defparam ram_block3a46.clk1_core_clock_enable = "ena1";
defparam ram_block3a46.data_interleave_offset_in_bits = 1;
defparam ram_block3a46.data_interleave_width_in_bits = 1;
defparam ram_block3a46.init_file = "meminit.hex";
defparam ram_block3a46.init_file_layout = "port_a";
defparam ram_block3a46.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a46.operation_mode = "bidir_dual_port";
defparam ram_block3a46.port_a_address_clear = "none";
defparam ram_block3a46.port_a_address_width = 13;
defparam ram_block3a46.port_a_byte_enable_clock = "none";
defparam ram_block3a46.port_a_data_out_clear = "none";
defparam ram_block3a46.port_a_data_out_clock = "none";
defparam ram_block3a46.port_a_data_width = 1;
defparam ram_block3a46.port_a_first_address = 0;
defparam ram_block3a46.port_a_first_bit_number = 14;
defparam ram_block3a46.port_a_last_address = 8191;
defparam ram_block3a46.port_a_logical_ram_depth = 16384;
defparam ram_block3a46.port_a_logical_ram_width = 32;
defparam ram_block3a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_address_clear = "none";
defparam ram_block3a46.port_b_address_clock = "clock1";
defparam ram_block3a46.port_b_address_width = 13;
defparam ram_block3a46.port_b_data_in_clock = "clock1";
defparam ram_block3a46.port_b_data_out_clear = "none";
defparam ram_block3a46.port_b_data_out_clock = "none";
defparam ram_block3a46.port_b_data_width = 1;
defparam ram_block3a46.port_b_first_address = 0;
defparam ram_block3a46.port_b_first_bit_number = 14;
defparam ram_block3a46.port_b_last_address = 8191;
defparam ram_block3a46.port_b_logical_ram_depth = 16384;
defparam ram_block3a46.port_b_logical_ram_width = 32;
defparam ram_block3a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_read_enable_clock = "clock1";
defparam ram_block3a46.port_b_write_enable_clock = "clock1";
defparam ram_block3a46.ram_block_type = "M9K";
defparam ram_block3a46.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y31_N0
cycloneive_ram_block ram_block3a14(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a14_PORTADATAOUT_bus),
	.portbdataout(ram_block3a14_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a14.clk0_core_clock_enable = "ena0";
defparam ram_block3a14.clk1_core_clock_enable = "ena1";
defparam ram_block3a14.data_interleave_offset_in_bits = 1;
defparam ram_block3a14.data_interleave_width_in_bits = 1;
defparam ram_block3a14.init_file = "meminit.hex";
defparam ram_block3a14.init_file_layout = "port_a";
defparam ram_block3a14.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a14.operation_mode = "bidir_dual_port";
defparam ram_block3a14.port_a_address_clear = "none";
defparam ram_block3a14.port_a_address_width = 13;
defparam ram_block3a14.port_a_byte_enable_clock = "none";
defparam ram_block3a14.port_a_data_out_clear = "none";
defparam ram_block3a14.port_a_data_out_clock = "none";
defparam ram_block3a14.port_a_data_width = 1;
defparam ram_block3a14.port_a_first_address = 0;
defparam ram_block3a14.port_a_first_bit_number = 14;
defparam ram_block3a14.port_a_last_address = 8191;
defparam ram_block3a14.port_a_logical_ram_depth = 16384;
defparam ram_block3a14.port_a_logical_ram_width = 32;
defparam ram_block3a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_address_clear = "none";
defparam ram_block3a14.port_b_address_clock = "clock1";
defparam ram_block3a14.port_b_address_width = 13;
defparam ram_block3a14.port_b_data_in_clock = "clock1";
defparam ram_block3a14.port_b_data_out_clear = "none";
defparam ram_block3a14.port_b_data_out_clock = "none";
defparam ram_block3a14.port_b_data_width = 1;
defparam ram_block3a14.port_b_first_address = 0;
defparam ram_block3a14.port_b_first_bit_number = 14;
defparam ram_block3a14.port_b_last_address = 8191;
defparam ram_block3a14.port_b_logical_ram_depth = 16384;
defparam ram_block3a14.port_b_logical_ram_width = 32;
defparam ram_block3a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_read_enable_clock = "clock1";
defparam ram_block3a14.port_b_write_enable_clock = "clock1";
defparam ram_block3a14.ram_block_type = "M9K";
defparam ram_block3a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000224A200503;
// synopsys translate_on

// Location: M9K_X78_Y30_N0
cycloneive_ram_block ram_block3a47(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a47_PORTADATAOUT_bus),
	.portbdataout(ram_block3a47_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a47.clk0_core_clock_enable = "ena0";
defparam ram_block3a47.clk1_core_clock_enable = "ena1";
defparam ram_block3a47.data_interleave_offset_in_bits = 1;
defparam ram_block3a47.data_interleave_width_in_bits = 1;
defparam ram_block3a47.init_file = "meminit.hex";
defparam ram_block3a47.init_file_layout = "port_a";
defparam ram_block3a47.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a47.operation_mode = "bidir_dual_port";
defparam ram_block3a47.port_a_address_clear = "none";
defparam ram_block3a47.port_a_address_width = 13;
defparam ram_block3a47.port_a_byte_enable_clock = "none";
defparam ram_block3a47.port_a_data_out_clear = "none";
defparam ram_block3a47.port_a_data_out_clock = "none";
defparam ram_block3a47.port_a_data_width = 1;
defparam ram_block3a47.port_a_first_address = 0;
defparam ram_block3a47.port_a_first_bit_number = 15;
defparam ram_block3a47.port_a_last_address = 8191;
defparam ram_block3a47.port_a_logical_ram_depth = 16384;
defparam ram_block3a47.port_a_logical_ram_width = 32;
defparam ram_block3a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_address_clear = "none";
defparam ram_block3a47.port_b_address_clock = "clock1";
defparam ram_block3a47.port_b_address_width = 13;
defparam ram_block3a47.port_b_data_in_clock = "clock1";
defparam ram_block3a47.port_b_data_out_clear = "none";
defparam ram_block3a47.port_b_data_out_clock = "none";
defparam ram_block3a47.port_b_data_width = 1;
defparam ram_block3a47.port_b_first_address = 0;
defparam ram_block3a47.port_b_first_bit_number = 15;
defparam ram_block3a47.port_b_last_address = 8191;
defparam ram_block3a47.port_b_logical_ram_depth = 16384;
defparam ram_block3a47.port_b_logical_ram_width = 32;
defparam ram_block3a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_read_enable_clock = "clock1";
defparam ram_block3a47.port_b_write_enable_clock = "clock1";
defparam ram_block3a47.ram_block_type = "M9K";
defparam ram_block3a47.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y31_N0
cycloneive_ram_block ram_block3a15(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a15_PORTADATAOUT_bus),
	.portbdataout(ram_block3a15_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a15.clk0_core_clock_enable = "ena0";
defparam ram_block3a15.clk1_core_clock_enable = "ena1";
defparam ram_block3a15.data_interleave_offset_in_bits = 1;
defparam ram_block3a15.data_interleave_width_in_bits = 1;
defparam ram_block3a15.init_file = "meminit.hex";
defparam ram_block3a15.init_file_layout = "port_a";
defparam ram_block3a15.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a15.operation_mode = "bidir_dual_port";
defparam ram_block3a15.port_a_address_clear = "none";
defparam ram_block3a15.port_a_address_width = 13;
defparam ram_block3a15.port_a_byte_enable_clock = "none";
defparam ram_block3a15.port_a_data_out_clear = "none";
defparam ram_block3a15.port_a_data_out_clock = "none";
defparam ram_block3a15.port_a_data_width = 1;
defparam ram_block3a15.port_a_first_address = 0;
defparam ram_block3a15.port_a_first_bit_number = 15;
defparam ram_block3a15.port_a_last_address = 8191;
defparam ram_block3a15.port_a_logical_ram_depth = 16384;
defparam ram_block3a15.port_a_logical_ram_width = 32;
defparam ram_block3a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_address_clear = "none";
defparam ram_block3a15.port_b_address_clock = "clock1";
defparam ram_block3a15.port_b_address_width = 13;
defparam ram_block3a15.port_b_data_in_clock = "clock1";
defparam ram_block3a15.port_b_data_out_clear = "none";
defparam ram_block3a15.port_b_data_out_clock = "none";
defparam ram_block3a15.port_b_data_width = 1;
defparam ram_block3a15.port_b_first_address = 0;
defparam ram_block3a15.port_b_first_bit_number = 15;
defparam ram_block3a15.port_b_last_address = 8191;
defparam ram_block3a15.port_b_logical_ram_depth = 16384;
defparam ram_block3a15.port_b_logical_ram_width = 32;
defparam ram_block3a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_read_enable_clock = "clock1";
defparam ram_block3a15.port_b_write_enable_clock = "clock1";
defparam ram_block3a15.ram_block_type = "M9K";
defparam ram_block3a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002042100002242206063;
// synopsys translate_on

// Location: M9K_X51_Y27_N0
cycloneive_ram_block ram_block3a48(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a48_PORTADATAOUT_bus),
	.portbdataout(ram_block3a48_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a48.clk0_core_clock_enable = "ena0";
defparam ram_block3a48.clk1_core_clock_enable = "ena1";
defparam ram_block3a48.data_interleave_offset_in_bits = 1;
defparam ram_block3a48.data_interleave_width_in_bits = 1;
defparam ram_block3a48.init_file = "meminit.hex";
defparam ram_block3a48.init_file_layout = "port_a";
defparam ram_block3a48.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a48.operation_mode = "bidir_dual_port";
defparam ram_block3a48.port_a_address_clear = "none";
defparam ram_block3a48.port_a_address_width = 13;
defparam ram_block3a48.port_a_byte_enable_clock = "none";
defparam ram_block3a48.port_a_data_out_clear = "none";
defparam ram_block3a48.port_a_data_out_clock = "none";
defparam ram_block3a48.port_a_data_width = 1;
defparam ram_block3a48.port_a_first_address = 0;
defparam ram_block3a48.port_a_first_bit_number = 16;
defparam ram_block3a48.port_a_last_address = 8191;
defparam ram_block3a48.port_a_logical_ram_depth = 16384;
defparam ram_block3a48.port_a_logical_ram_width = 32;
defparam ram_block3a48.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_address_clear = "none";
defparam ram_block3a48.port_b_address_clock = "clock1";
defparam ram_block3a48.port_b_address_width = 13;
defparam ram_block3a48.port_b_data_in_clock = "clock1";
defparam ram_block3a48.port_b_data_out_clear = "none";
defparam ram_block3a48.port_b_data_out_clock = "none";
defparam ram_block3a48.port_b_data_width = 1;
defparam ram_block3a48.port_b_first_address = 0;
defparam ram_block3a48.port_b_first_bit_number = 16;
defparam ram_block3a48.port_b_last_address = 8191;
defparam ram_block3a48.port_b_logical_ram_depth = 16384;
defparam ram_block3a48.port_b_logical_ram_width = 32;
defparam ram_block3a48.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_read_enable_clock = "clock1";
defparam ram_block3a48.port_b_write_enable_clock = "clock1";
defparam ram_block3a48.ram_block_type = "M9K";
defparam ram_block3a48.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y25_N0
cycloneive_ram_block ram_block3a16(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a16_PORTADATAOUT_bus),
	.portbdataout(ram_block3a16_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a16.clk0_core_clock_enable = "ena0";
defparam ram_block3a16.clk1_core_clock_enable = "ena1";
defparam ram_block3a16.data_interleave_offset_in_bits = 1;
defparam ram_block3a16.data_interleave_width_in_bits = 1;
defparam ram_block3a16.init_file = "meminit.hex";
defparam ram_block3a16.init_file_layout = "port_a";
defparam ram_block3a16.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a16.operation_mode = "bidir_dual_port";
defparam ram_block3a16.port_a_address_clear = "none";
defparam ram_block3a16.port_a_address_width = 13;
defparam ram_block3a16.port_a_byte_enable_clock = "none";
defparam ram_block3a16.port_a_data_out_clear = "none";
defparam ram_block3a16.port_a_data_out_clock = "none";
defparam ram_block3a16.port_a_data_width = 1;
defparam ram_block3a16.port_a_first_address = 0;
defparam ram_block3a16.port_a_first_bit_number = 16;
defparam ram_block3a16.port_a_last_address = 8191;
defparam ram_block3a16.port_a_logical_ram_depth = 16384;
defparam ram_block3a16.port_a_logical_ram_width = 32;
defparam ram_block3a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_address_clear = "none";
defparam ram_block3a16.port_b_address_clock = "clock1";
defparam ram_block3a16.port_b_address_width = 13;
defparam ram_block3a16.port_b_data_in_clock = "clock1";
defparam ram_block3a16.port_b_data_out_clear = "none";
defparam ram_block3a16.port_b_data_out_clock = "none";
defparam ram_block3a16.port_b_data_width = 1;
defparam ram_block3a16.port_b_first_address = 0;
defparam ram_block3a16.port_b_first_bit_number = 16;
defparam ram_block3a16.port_b_last_address = 8191;
defparam ram_block3a16.port_b_logical_ram_depth = 16384;
defparam ram_block3a16.port_b_logical_ram_width = 32;
defparam ram_block3a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_read_enable_clock = "clock1";
defparam ram_block3a16.port_b_write_enable_clock = "clock1";
defparam ram_block3a16.ram_block_type = "M9K";
defparam ram_block3a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000205A122003613254042;
// synopsys translate_on

// Location: M9K_X51_Y28_N0
cycloneive_ram_block ram_block3a49(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a49_PORTADATAOUT_bus),
	.portbdataout(ram_block3a49_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a49.clk0_core_clock_enable = "ena0";
defparam ram_block3a49.clk1_core_clock_enable = "ena1";
defparam ram_block3a49.data_interleave_offset_in_bits = 1;
defparam ram_block3a49.data_interleave_width_in_bits = 1;
defparam ram_block3a49.init_file = "meminit.hex";
defparam ram_block3a49.init_file_layout = "port_a";
defparam ram_block3a49.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a49.operation_mode = "bidir_dual_port";
defparam ram_block3a49.port_a_address_clear = "none";
defparam ram_block3a49.port_a_address_width = 13;
defparam ram_block3a49.port_a_byte_enable_clock = "none";
defparam ram_block3a49.port_a_data_out_clear = "none";
defparam ram_block3a49.port_a_data_out_clock = "none";
defparam ram_block3a49.port_a_data_width = 1;
defparam ram_block3a49.port_a_first_address = 0;
defparam ram_block3a49.port_a_first_bit_number = 17;
defparam ram_block3a49.port_a_last_address = 8191;
defparam ram_block3a49.port_a_logical_ram_depth = 16384;
defparam ram_block3a49.port_a_logical_ram_width = 32;
defparam ram_block3a49.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_address_clear = "none";
defparam ram_block3a49.port_b_address_clock = "clock1";
defparam ram_block3a49.port_b_address_width = 13;
defparam ram_block3a49.port_b_data_in_clock = "clock1";
defparam ram_block3a49.port_b_data_out_clear = "none";
defparam ram_block3a49.port_b_data_out_clock = "none";
defparam ram_block3a49.port_b_data_width = 1;
defparam ram_block3a49.port_b_first_address = 0;
defparam ram_block3a49.port_b_first_bit_number = 17;
defparam ram_block3a49.port_b_last_address = 8191;
defparam ram_block3a49.port_b_logical_ram_depth = 16384;
defparam ram_block3a49.port_b_logical_ram_width = 32;
defparam ram_block3a49.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_read_enable_clock = "clock1";
defparam ram_block3a49.port_b_write_enable_clock = "clock1";
defparam ram_block3a49.ram_block_type = "M9K";
defparam ram_block3a49.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y26_N0
cycloneive_ram_block ram_block3a17(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a17_PORTADATAOUT_bus),
	.portbdataout(ram_block3a17_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a17.clk0_core_clock_enable = "ena0";
defparam ram_block3a17.clk1_core_clock_enable = "ena1";
defparam ram_block3a17.data_interleave_offset_in_bits = 1;
defparam ram_block3a17.data_interleave_width_in_bits = 1;
defparam ram_block3a17.init_file = "meminit.hex";
defparam ram_block3a17.init_file_layout = "port_a";
defparam ram_block3a17.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a17.operation_mode = "bidir_dual_port";
defparam ram_block3a17.port_a_address_clear = "none";
defparam ram_block3a17.port_a_address_width = 13;
defparam ram_block3a17.port_a_byte_enable_clock = "none";
defparam ram_block3a17.port_a_data_out_clear = "none";
defparam ram_block3a17.port_a_data_out_clock = "none";
defparam ram_block3a17.port_a_data_width = 1;
defparam ram_block3a17.port_a_first_address = 0;
defparam ram_block3a17.port_a_first_bit_number = 17;
defparam ram_block3a17.port_a_last_address = 8191;
defparam ram_block3a17.port_a_logical_ram_depth = 16384;
defparam ram_block3a17.port_a_logical_ram_width = 32;
defparam ram_block3a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_address_clear = "none";
defparam ram_block3a17.port_b_address_clock = "clock1";
defparam ram_block3a17.port_b_address_width = 13;
defparam ram_block3a17.port_b_data_in_clock = "clock1";
defparam ram_block3a17.port_b_data_out_clear = "none";
defparam ram_block3a17.port_b_data_out_clock = "none";
defparam ram_block3a17.port_b_data_width = 1;
defparam ram_block3a17.port_b_first_address = 0;
defparam ram_block3a17.port_b_first_bit_number = 17;
defparam ram_block3a17.port_b_last_address = 8191;
defparam ram_block3a17.port_b_logical_ram_depth = 16384;
defparam ram_block3a17.port_b_logical_ram_width = 32;
defparam ram_block3a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_read_enable_clock = "clock1";
defparam ram_block3a17.port_b_write_enable_clock = "clock1";
defparam ram_block3a17.ram_block_type = "M9K";
defparam ram_block3a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006C0340C001602060001;
// synopsys translate_on

// Location: M9K_X78_Y39_N0
cycloneive_ram_block ram_block3a50(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a50_PORTADATAOUT_bus),
	.portbdataout(ram_block3a50_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a50.clk0_core_clock_enable = "ena0";
defparam ram_block3a50.clk1_core_clock_enable = "ena1";
defparam ram_block3a50.data_interleave_offset_in_bits = 1;
defparam ram_block3a50.data_interleave_width_in_bits = 1;
defparam ram_block3a50.init_file = "meminit.hex";
defparam ram_block3a50.init_file_layout = "port_a";
defparam ram_block3a50.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a50.operation_mode = "bidir_dual_port";
defparam ram_block3a50.port_a_address_clear = "none";
defparam ram_block3a50.port_a_address_width = 13;
defparam ram_block3a50.port_a_byte_enable_clock = "none";
defparam ram_block3a50.port_a_data_out_clear = "none";
defparam ram_block3a50.port_a_data_out_clock = "none";
defparam ram_block3a50.port_a_data_width = 1;
defparam ram_block3a50.port_a_first_address = 0;
defparam ram_block3a50.port_a_first_bit_number = 18;
defparam ram_block3a50.port_a_last_address = 8191;
defparam ram_block3a50.port_a_logical_ram_depth = 16384;
defparam ram_block3a50.port_a_logical_ram_width = 32;
defparam ram_block3a50.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_address_clear = "none";
defparam ram_block3a50.port_b_address_clock = "clock1";
defparam ram_block3a50.port_b_address_width = 13;
defparam ram_block3a50.port_b_data_in_clock = "clock1";
defparam ram_block3a50.port_b_data_out_clear = "none";
defparam ram_block3a50.port_b_data_out_clock = "none";
defparam ram_block3a50.port_b_data_width = 1;
defparam ram_block3a50.port_b_first_address = 0;
defparam ram_block3a50.port_b_first_bit_number = 18;
defparam ram_block3a50.port_b_last_address = 8191;
defparam ram_block3a50.port_b_logical_ram_depth = 16384;
defparam ram_block3a50.port_b_logical_ram_width = 32;
defparam ram_block3a50.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_read_enable_clock = "clock1";
defparam ram_block3a50.port_b_write_enable_clock = "clock1";
defparam ram_block3a50.ram_block_type = "M9K";
defparam ram_block3a50.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y41_N0
cycloneive_ram_block ram_block3a18(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a18_PORTADATAOUT_bus),
	.portbdataout(ram_block3a18_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a18.clk0_core_clock_enable = "ena0";
defparam ram_block3a18.clk1_core_clock_enable = "ena1";
defparam ram_block3a18.data_interleave_offset_in_bits = 1;
defparam ram_block3a18.data_interleave_width_in_bits = 1;
defparam ram_block3a18.init_file = "meminit.hex";
defparam ram_block3a18.init_file_layout = "port_a";
defparam ram_block3a18.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a18.operation_mode = "bidir_dual_port";
defparam ram_block3a18.port_a_address_clear = "none";
defparam ram_block3a18.port_a_address_width = 13;
defparam ram_block3a18.port_a_byte_enable_clock = "none";
defparam ram_block3a18.port_a_data_out_clear = "none";
defparam ram_block3a18.port_a_data_out_clock = "none";
defparam ram_block3a18.port_a_data_width = 1;
defparam ram_block3a18.port_a_first_address = 0;
defparam ram_block3a18.port_a_first_bit_number = 18;
defparam ram_block3a18.port_a_last_address = 8191;
defparam ram_block3a18.port_a_logical_ram_depth = 16384;
defparam ram_block3a18.port_a_logical_ram_width = 32;
defparam ram_block3a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_address_clear = "none";
defparam ram_block3a18.port_b_address_clock = "clock1";
defparam ram_block3a18.port_b_address_width = 13;
defparam ram_block3a18.port_b_data_in_clock = "clock1";
defparam ram_block3a18.port_b_data_out_clear = "none";
defparam ram_block3a18.port_b_data_out_clock = "none";
defparam ram_block3a18.port_b_data_width = 1;
defparam ram_block3a18.port_b_first_address = 0;
defparam ram_block3a18.port_b_first_bit_number = 18;
defparam ram_block3a18.port_b_last_address = 8191;
defparam ram_block3a18.port_b_logical_ram_depth = 16384;
defparam ram_block3a18.port_b_logical_ram_width = 32;
defparam ram_block3a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_read_enable_clock = "clock1";
defparam ram_block3a18.port_b_write_enable_clock = "clock1";
defparam ram_block3a18.ram_block_type = "M9K";
defparam ram_block3a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060C3180001703286867;
// synopsys translate_on

// Location: M9K_X78_Y36_N0
cycloneive_ram_block ram_block3a51(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a51_PORTADATAOUT_bus),
	.portbdataout(ram_block3a51_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a51.clk0_core_clock_enable = "ena0";
defparam ram_block3a51.clk1_core_clock_enable = "ena1";
defparam ram_block3a51.data_interleave_offset_in_bits = 1;
defparam ram_block3a51.data_interleave_width_in_bits = 1;
defparam ram_block3a51.init_file = "meminit.hex";
defparam ram_block3a51.init_file_layout = "port_a";
defparam ram_block3a51.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a51.operation_mode = "bidir_dual_port";
defparam ram_block3a51.port_a_address_clear = "none";
defparam ram_block3a51.port_a_address_width = 13;
defparam ram_block3a51.port_a_byte_enable_clock = "none";
defparam ram_block3a51.port_a_data_out_clear = "none";
defparam ram_block3a51.port_a_data_out_clock = "none";
defparam ram_block3a51.port_a_data_width = 1;
defparam ram_block3a51.port_a_first_address = 0;
defparam ram_block3a51.port_a_first_bit_number = 19;
defparam ram_block3a51.port_a_last_address = 8191;
defparam ram_block3a51.port_a_logical_ram_depth = 16384;
defparam ram_block3a51.port_a_logical_ram_width = 32;
defparam ram_block3a51.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_address_clear = "none";
defparam ram_block3a51.port_b_address_clock = "clock1";
defparam ram_block3a51.port_b_address_width = 13;
defparam ram_block3a51.port_b_data_in_clock = "clock1";
defparam ram_block3a51.port_b_data_out_clear = "none";
defparam ram_block3a51.port_b_data_out_clock = "none";
defparam ram_block3a51.port_b_data_width = 1;
defparam ram_block3a51.port_b_first_address = 0;
defparam ram_block3a51.port_b_first_bit_number = 19;
defparam ram_block3a51.port_b_last_address = 8191;
defparam ram_block3a51.port_b_logical_ram_depth = 16384;
defparam ram_block3a51.port_b_logical_ram_width = 32;
defparam ram_block3a51.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_read_enable_clock = "clock1";
defparam ram_block3a51.port_b_write_enable_clock = "clock1";
defparam ram_block3a51.ram_block_type = "M9K";
defparam ram_block3a51.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y35_N0
cycloneive_ram_block ram_block3a19(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a19_PORTADATAOUT_bus),
	.portbdataout(ram_block3a19_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a19.clk0_core_clock_enable = "ena0";
defparam ram_block3a19.clk1_core_clock_enable = "ena1";
defparam ram_block3a19.data_interleave_offset_in_bits = 1;
defparam ram_block3a19.data_interleave_width_in_bits = 1;
defparam ram_block3a19.init_file = "meminit.hex";
defparam ram_block3a19.init_file_layout = "port_a";
defparam ram_block3a19.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a19.operation_mode = "bidir_dual_port";
defparam ram_block3a19.port_a_address_clear = "none";
defparam ram_block3a19.port_a_address_width = 13;
defparam ram_block3a19.port_a_byte_enable_clock = "none";
defparam ram_block3a19.port_a_data_out_clear = "none";
defparam ram_block3a19.port_a_data_out_clock = "none";
defparam ram_block3a19.port_a_data_width = 1;
defparam ram_block3a19.port_a_first_address = 0;
defparam ram_block3a19.port_a_first_bit_number = 19;
defparam ram_block3a19.port_a_last_address = 8191;
defparam ram_block3a19.port_a_logical_ram_depth = 16384;
defparam ram_block3a19.port_a_logical_ram_width = 32;
defparam ram_block3a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_address_clear = "none";
defparam ram_block3a19.port_b_address_clock = "clock1";
defparam ram_block3a19.port_b_address_width = 13;
defparam ram_block3a19.port_b_data_in_clock = "clock1";
defparam ram_block3a19.port_b_data_out_clear = "none";
defparam ram_block3a19.port_b_data_out_clock = "none";
defparam ram_block3a19.port_b_data_width = 1;
defparam ram_block3a19.port_b_first_address = 0;
defparam ram_block3a19.port_b_first_bit_number = 19;
defparam ram_block3a19.port_b_last_address = 8191;
defparam ram_block3a19.port_b_logical_ram_depth = 16384;
defparam ram_block3a19.port_b_logical_ram_width = 32;
defparam ram_block3a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_read_enable_clock = "clock1";
defparam ram_block3a19.port_b_write_enable_clock = "clock1";
defparam ram_block3a19.ram_block_type = "M9K";
defparam ram_block3a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001C38C6E09B6D7701203;
// synopsys translate_on

// Location: M9K_X51_Y37_N0
cycloneive_ram_block ram_block3a52(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a52_PORTADATAOUT_bus),
	.portbdataout(ram_block3a52_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a52.clk0_core_clock_enable = "ena0";
defparam ram_block3a52.clk1_core_clock_enable = "ena1";
defparam ram_block3a52.data_interleave_offset_in_bits = 1;
defparam ram_block3a52.data_interleave_width_in_bits = 1;
defparam ram_block3a52.init_file = "meminit.hex";
defparam ram_block3a52.init_file_layout = "port_a";
defparam ram_block3a52.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a52.operation_mode = "bidir_dual_port";
defparam ram_block3a52.port_a_address_clear = "none";
defparam ram_block3a52.port_a_address_width = 13;
defparam ram_block3a52.port_a_byte_enable_clock = "none";
defparam ram_block3a52.port_a_data_out_clear = "none";
defparam ram_block3a52.port_a_data_out_clock = "none";
defparam ram_block3a52.port_a_data_width = 1;
defparam ram_block3a52.port_a_first_address = 0;
defparam ram_block3a52.port_a_first_bit_number = 20;
defparam ram_block3a52.port_a_last_address = 8191;
defparam ram_block3a52.port_a_logical_ram_depth = 16384;
defparam ram_block3a52.port_a_logical_ram_width = 32;
defparam ram_block3a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_address_clear = "none";
defparam ram_block3a52.port_b_address_clock = "clock1";
defparam ram_block3a52.port_b_address_width = 13;
defparam ram_block3a52.port_b_data_in_clock = "clock1";
defparam ram_block3a52.port_b_data_out_clear = "none";
defparam ram_block3a52.port_b_data_out_clock = "none";
defparam ram_block3a52.port_b_data_width = 1;
defparam ram_block3a52.port_b_first_address = 0;
defparam ram_block3a52.port_b_first_bit_number = 20;
defparam ram_block3a52.port_b_last_address = 8191;
defparam ram_block3a52.port_b_logical_ram_depth = 16384;
defparam ram_block3a52.port_b_logical_ram_width = 32;
defparam ram_block3a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_read_enable_clock = "clock1";
defparam ram_block3a52.port_b_write_enable_clock = "clock1";
defparam ram_block3a52.ram_block_type = "M9K";
defparam ram_block3a52.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y39_N0
cycloneive_ram_block ram_block3a20(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a20_PORTADATAOUT_bus),
	.portbdataout(ram_block3a20_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a20.clk0_core_clock_enable = "ena0";
defparam ram_block3a20.clk1_core_clock_enable = "ena1";
defparam ram_block3a20.data_interleave_offset_in_bits = 1;
defparam ram_block3a20.data_interleave_width_in_bits = 1;
defparam ram_block3a20.init_file = "meminit.hex";
defparam ram_block3a20.init_file_layout = "port_a";
defparam ram_block3a20.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a20.operation_mode = "bidir_dual_port";
defparam ram_block3a20.port_a_address_clear = "none";
defparam ram_block3a20.port_a_address_width = 13;
defparam ram_block3a20.port_a_byte_enable_clock = "none";
defparam ram_block3a20.port_a_data_out_clear = "none";
defparam ram_block3a20.port_a_data_out_clock = "none";
defparam ram_block3a20.port_a_data_width = 1;
defparam ram_block3a20.port_a_first_address = 0;
defparam ram_block3a20.port_a_first_bit_number = 20;
defparam ram_block3a20.port_a_last_address = 8191;
defparam ram_block3a20.port_a_logical_ram_depth = 16384;
defparam ram_block3a20.port_a_logical_ram_width = 32;
defparam ram_block3a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_address_clear = "none";
defparam ram_block3a20.port_b_address_clock = "clock1";
defparam ram_block3a20.port_b_address_width = 13;
defparam ram_block3a20.port_b_data_in_clock = "clock1";
defparam ram_block3a20.port_b_data_out_clear = "none";
defparam ram_block3a20.port_b_data_out_clock = "none";
defparam ram_block3a20.port_b_data_width = 1;
defparam ram_block3a20.port_b_first_address = 0;
defparam ram_block3a20.port_b_first_bit_number = 20;
defparam ram_block3a20.port_b_last_address = 8191;
defparam ram_block3a20.port_b_logical_ram_depth = 16384;
defparam ram_block3a20.port_b_logical_ram_width = 32;
defparam ram_block3a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_read_enable_clock = "clock1";
defparam ram_block3a20.port_b_write_enable_clock = "clock1";
defparam ram_block3a20.ram_block_type = "M9K";
defparam ram_block3a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A0832F000B;
// synopsys translate_on

// Location: M9K_X51_Y36_N0
cycloneive_ram_block ram_block3a53(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a53_PORTADATAOUT_bus),
	.portbdataout(ram_block3a53_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a53.clk0_core_clock_enable = "ena0";
defparam ram_block3a53.clk1_core_clock_enable = "ena1";
defparam ram_block3a53.data_interleave_offset_in_bits = 1;
defparam ram_block3a53.data_interleave_width_in_bits = 1;
defparam ram_block3a53.init_file = "meminit.hex";
defparam ram_block3a53.init_file_layout = "port_a";
defparam ram_block3a53.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a53.operation_mode = "bidir_dual_port";
defparam ram_block3a53.port_a_address_clear = "none";
defparam ram_block3a53.port_a_address_width = 13;
defparam ram_block3a53.port_a_byte_enable_clock = "none";
defparam ram_block3a53.port_a_data_out_clear = "none";
defparam ram_block3a53.port_a_data_out_clock = "none";
defparam ram_block3a53.port_a_data_width = 1;
defparam ram_block3a53.port_a_first_address = 0;
defparam ram_block3a53.port_a_first_bit_number = 21;
defparam ram_block3a53.port_a_last_address = 8191;
defparam ram_block3a53.port_a_logical_ram_depth = 16384;
defparam ram_block3a53.port_a_logical_ram_width = 32;
defparam ram_block3a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_address_clear = "none";
defparam ram_block3a53.port_b_address_clock = "clock1";
defparam ram_block3a53.port_b_address_width = 13;
defparam ram_block3a53.port_b_data_in_clock = "clock1";
defparam ram_block3a53.port_b_data_out_clear = "none";
defparam ram_block3a53.port_b_data_out_clock = "none";
defparam ram_block3a53.port_b_data_width = 1;
defparam ram_block3a53.port_b_first_address = 0;
defparam ram_block3a53.port_b_first_bit_number = 21;
defparam ram_block3a53.port_b_last_address = 8191;
defparam ram_block3a53.port_b_logical_ram_depth = 16384;
defparam ram_block3a53.port_b_logical_ram_width = 32;
defparam ram_block3a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_read_enable_clock = "clock1";
defparam ram_block3a53.port_b_write_enable_clock = "clock1";
defparam ram_block3a53.ram_block_type = "M9K";
defparam ram_block3a53.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y35_N0
cycloneive_ram_block ram_block3a21(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a21_PORTADATAOUT_bus),
	.portbdataout(ram_block3a21_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a21.clk0_core_clock_enable = "ena0";
defparam ram_block3a21.clk1_core_clock_enable = "ena1";
defparam ram_block3a21.data_interleave_offset_in_bits = 1;
defparam ram_block3a21.data_interleave_width_in_bits = 1;
defparam ram_block3a21.init_file = "meminit.hex";
defparam ram_block3a21.init_file_layout = "port_a";
defparam ram_block3a21.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a21.operation_mode = "bidir_dual_port";
defparam ram_block3a21.port_a_address_clear = "none";
defparam ram_block3a21.port_a_address_width = 13;
defparam ram_block3a21.port_a_byte_enable_clock = "none";
defparam ram_block3a21.port_a_data_out_clear = "none";
defparam ram_block3a21.port_a_data_out_clock = "none";
defparam ram_block3a21.port_a_data_width = 1;
defparam ram_block3a21.port_a_first_address = 0;
defparam ram_block3a21.port_a_first_bit_number = 21;
defparam ram_block3a21.port_a_last_address = 8191;
defparam ram_block3a21.port_a_logical_ram_depth = 16384;
defparam ram_block3a21.port_a_logical_ram_width = 32;
defparam ram_block3a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_address_clear = "none";
defparam ram_block3a21.port_b_address_clock = "clock1";
defparam ram_block3a21.port_b_address_width = 13;
defparam ram_block3a21.port_b_data_in_clock = "clock1";
defparam ram_block3a21.port_b_data_out_clear = "none";
defparam ram_block3a21.port_b_data_out_clock = "none";
defparam ram_block3a21.port_b_data_width = 1;
defparam ram_block3a21.port_b_first_address = 0;
defparam ram_block3a21.port_b_first_bit_number = 21;
defparam ram_block3a21.port_b_last_address = 8191;
defparam ram_block3a21.port_b_logical_ram_depth = 16384;
defparam ram_block3a21.port_b_logical_ram_width = 32;
defparam ram_block3a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_read_enable_clock = "clock1";
defparam ram_block3a21.port_b_write_enable_clock = "clock1";
defparam ram_block3a21.ram_block_type = "M9K";
defparam ram_block3a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002A142119BCBBAB600000;
// synopsys translate_on

// Location: M9K_X64_Y33_N0
cycloneive_ram_block ram_block3a54(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a54_PORTADATAOUT_bus),
	.portbdataout(ram_block3a54_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a54.clk0_core_clock_enable = "ena0";
defparam ram_block3a54.clk1_core_clock_enable = "ena1";
defparam ram_block3a54.data_interleave_offset_in_bits = 1;
defparam ram_block3a54.data_interleave_width_in_bits = 1;
defparam ram_block3a54.init_file = "meminit.hex";
defparam ram_block3a54.init_file_layout = "port_a";
defparam ram_block3a54.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a54.operation_mode = "bidir_dual_port";
defparam ram_block3a54.port_a_address_clear = "none";
defparam ram_block3a54.port_a_address_width = 13;
defparam ram_block3a54.port_a_byte_enable_clock = "none";
defparam ram_block3a54.port_a_data_out_clear = "none";
defparam ram_block3a54.port_a_data_out_clock = "none";
defparam ram_block3a54.port_a_data_width = 1;
defparam ram_block3a54.port_a_first_address = 0;
defparam ram_block3a54.port_a_first_bit_number = 22;
defparam ram_block3a54.port_a_last_address = 8191;
defparam ram_block3a54.port_a_logical_ram_depth = 16384;
defparam ram_block3a54.port_a_logical_ram_width = 32;
defparam ram_block3a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_address_clear = "none";
defparam ram_block3a54.port_b_address_clock = "clock1";
defparam ram_block3a54.port_b_address_width = 13;
defparam ram_block3a54.port_b_data_in_clock = "clock1";
defparam ram_block3a54.port_b_data_out_clear = "none";
defparam ram_block3a54.port_b_data_out_clock = "none";
defparam ram_block3a54.port_b_data_width = 1;
defparam ram_block3a54.port_b_first_address = 0;
defparam ram_block3a54.port_b_first_bit_number = 22;
defparam ram_block3a54.port_b_last_address = 8191;
defparam ram_block3a54.port_b_logical_ram_depth = 16384;
defparam ram_block3a54.port_b_logical_ram_width = 32;
defparam ram_block3a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_read_enable_clock = "clock1";
defparam ram_block3a54.port_b_write_enable_clock = "clock1";
defparam ram_block3a54.ram_block_type = "M9K";
defparam ram_block3a54.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y33_N0
cycloneive_ram_block ram_block3a22(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a22_PORTADATAOUT_bus),
	.portbdataout(ram_block3a22_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a22.clk0_core_clock_enable = "ena0";
defparam ram_block3a22.clk1_core_clock_enable = "ena1";
defparam ram_block3a22.data_interleave_offset_in_bits = 1;
defparam ram_block3a22.data_interleave_width_in_bits = 1;
defparam ram_block3a22.init_file = "meminit.hex";
defparam ram_block3a22.init_file_layout = "port_a";
defparam ram_block3a22.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a22.operation_mode = "bidir_dual_port";
defparam ram_block3a22.port_a_address_clear = "none";
defparam ram_block3a22.port_a_address_width = 13;
defparam ram_block3a22.port_a_byte_enable_clock = "none";
defparam ram_block3a22.port_a_data_out_clear = "none";
defparam ram_block3a22.port_a_data_out_clock = "none";
defparam ram_block3a22.port_a_data_width = 1;
defparam ram_block3a22.port_a_first_address = 0;
defparam ram_block3a22.port_a_first_bit_number = 22;
defparam ram_block3a22.port_a_last_address = 8191;
defparam ram_block3a22.port_a_logical_ram_depth = 16384;
defparam ram_block3a22.port_a_logical_ram_width = 32;
defparam ram_block3a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_address_clear = "none";
defparam ram_block3a22.port_b_address_clock = "clock1";
defparam ram_block3a22.port_b_address_width = 13;
defparam ram_block3a22.port_b_data_in_clock = "clock1";
defparam ram_block3a22.port_b_data_out_clear = "none";
defparam ram_block3a22.port_b_data_out_clock = "none";
defparam ram_block3a22.port_b_data_width = 1;
defparam ram_block3a22.port_b_first_address = 0;
defparam ram_block3a22.port_b_first_bit_number = 22;
defparam ram_block3a22.port_b_last_address = 8191;
defparam ram_block3a22.port_b_logical_ram_depth = 16384;
defparam ram_block3a22.port_b_logical_ram_width = 32;
defparam ram_block3a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_read_enable_clock = "clock1";
defparam ram_block3a22.port_b_write_enable_clock = "clock1";
defparam ram_block3a22.ram_block_type = "M9K";
defparam ram_block3a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002E403004A40002000000;
// synopsys translate_on

// Location: M9K_X51_Y29_N0
cycloneive_ram_block ram_block3a55(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a55_PORTADATAOUT_bus),
	.portbdataout(ram_block3a55_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a55.clk0_core_clock_enable = "ena0";
defparam ram_block3a55.clk1_core_clock_enable = "ena1";
defparam ram_block3a55.data_interleave_offset_in_bits = 1;
defparam ram_block3a55.data_interleave_width_in_bits = 1;
defparam ram_block3a55.init_file = "meminit.hex";
defparam ram_block3a55.init_file_layout = "port_a";
defparam ram_block3a55.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a55.operation_mode = "bidir_dual_port";
defparam ram_block3a55.port_a_address_clear = "none";
defparam ram_block3a55.port_a_address_width = 13;
defparam ram_block3a55.port_a_byte_enable_clock = "none";
defparam ram_block3a55.port_a_data_out_clear = "none";
defparam ram_block3a55.port_a_data_out_clock = "none";
defparam ram_block3a55.port_a_data_width = 1;
defparam ram_block3a55.port_a_first_address = 0;
defparam ram_block3a55.port_a_first_bit_number = 23;
defparam ram_block3a55.port_a_last_address = 8191;
defparam ram_block3a55.port_a_logical_ram_depth = 16384;
defparam ram_block3a55.port_a_logical_ram_width = 32;
defparam ram_block3a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_address_clear = "none";
defparam ram_block3a55.port_b_address_clock = "clock1";
defparam ram_block3a55.port_b_address_width = 13;
defparam ram_block3a55.port_b_data_in_clock = "clock1";
defparam ram_block3a55.port_b_data_out_clear = "none";
defparam ram_block3a55.port_b_data_out_clock = "none";
defparam ram_block3a55.port_b_data_width = 1;
defparam ram_block3a55.port_b_first_address = 0;
defparam ram_block3a55.port_b_first_bit_number = 23;
defparam ram_block3a55.port_b_last_address = 8191;
defparam ram_block3a55.port_b_logical_ram_depth = 16384;
defparam ram_block3a55.port_b_logical_ram_width = 32;
defparam ram_block3a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_read_enable_clock = "clock1";
defparam ram_block3a55.port_b_write_enable_clock = "clock1";
defparam ram_block3a55.ram_block_type = "M9K";
defparam ram_block3a55.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y29_N0
cycloneive_ram_block ram_block3a23(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a23_PORTADATAOUT_bus),
	.portbdataout(ram_block3a23_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a23.clk0_core_clock_enable = "ena0";
defparam ram_block3a23.clk1_core_clock_enable = "ena1";
defparam ram_block3a23.data_interleave_offset_in_bits = 1;
defparam ram_block3a23.data_interleave_width_in_bits = 1;
defparam ram_block3a23.init_file = "meminit.hex";
defparam ram_block3a23.init_file_layout = "port_a";
defparam ram_block3a23.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a23.operation_mode = "bidir_dual_port";
defparam ram_block3a23.port_a_address_clear = "none";
defparam ram_block3a23.port_a_address_width = 13;
defparam ram_block3a23.port_a_byte_enable_clock = "none";
defparam ram_block3a23.port_a_data_out_clear = "none";
defparam ram_block3a23.port_a_data_out_clock = "none";
defparam ram_block3a23.port_a_data_width = 1;
defparam ram_block3a23.port_a_first_address = 0;
defparam ram_block3a23.port_a_first_bit_number = 23;
defparam ram_block3a23.port_a_last_address = 8191;
defparam ram_block3a23.port_a_logical_ram_depth = 16384;
defparam ram_block3a23.port_a_logical_ram_width = 32;
defparam ram_block3a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_address_clear = "none";
defparam ram_block3a23.port_b_address_clock = "clock1";
defparam ram_block3a23.port_b_address_width = 13;
defparam ram_block3a23.port_b_data_in_clock = "clock1";
defparam ram_block3a23.port_b_data_out_clear = "none";
defparam ram_block3a23.port_b_data_out_clock = "none";
defparam ram_block3a23.port_b_data_width = 1;
defparam ram_block3a23.port_b_first_address = 0;
defparam ram_block3a23.port_b_first_bit_number = 23;
defparam ram_block3a23.port_b_last_address = 8191;
defparam ram_block3a23.port_b_logical_ram_depth = 16384;
defparam ram_block3a23.port_b_logical_ram_width = 32;
defparam ram_block3a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_read_enable_clock = "clock1";
defparam ram_block3a23.port_b_write_enable_clock = "clock1";
defparam ram_block3a23.ram_block_type = "M9K";
defparam ram_block3a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002E5CB187BC004B601000;
// synopsys translate_on

// Location: M9K_X64_Y37_N0
cycloneive_ram_block ram_block3a56(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a56_PORTADATAOUT_bus),
	.portbdataout(ram_block3a56_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a56.clk0_core_clock_enable = "ena0";
defparam ram_block3a56.clk1_core_clock_enable = "ena1";
defparam ram_block3a56.data_interleave_offset_in_bits = 1;
defparam ram_block3a56.data_interleave_width_in_bits = 1;
defparam ram_block3a56.init_file = "meminit.hex";
defparam ram_block3a56.init_file_layout = "port_a";
defparam ram_block3a56.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a56.operation_mode = "bidir_dual_port";
defparam ram_block3a56.port_a_address_clear = "none";
defparam ram_block3a56.port_a_address_width = 13;
defparam ram_block3a56.port_a_byte_enable_clock = "none";
defparam ram_block3a56.port_a_data_out_clear = "none";
defparam ram_block3a56.port_a_data_out_clock = "none";
defparam ram_block3a56.port_a_data_width = 1;
defparam ram_block3a56.port_a_first_address = 0;
defparam ram_block3a56.port_a_first_bit_number = 24;
defparam ram_block3a56.port_a_last_address = 8191;
defparam ram_block3a56.port_a_logical_ram_depth = 16384;
defparam ram_block3a56.port_a_logical_ram_width = 32;
defparam ram_block3a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_address_clear = "none";
defparam ram_block3a56.port_b_address_clock = "clock1";
defparam ram_block3a56.port_b_address_width = 13;
defparam ram_block3a56.port_b_data_in_clock = "clock1";
defparam ram_block3a56.port_b_data_out_clear = "none";
defparam ram_block3a56.port_b_data_out_clock = "none";
defparam ram_block3a56.port_b_data_width = 1;
defparam ram_block3a56.port_b_first_address = 0;
defparam ram_block3a56.port_b_first_bit_number = 24;
defparam ram_block3a56.port_b_last_address = 8191;
defparam ram_block3a56.port_b_logical_ram_depth = 16384;
defparam ram_block3a56.port_b_logical_ram_width = 32;
defparam ram_block3a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_read_enable_clock = "clock1";
defparam ram_block3a56.port_b_write_enable_clock = "clock1";
defparam ram_block3a56.ram_block_type = "M9K";
defparam ram_block3a56.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y37_N0
cycloneive_ram_block ram_block3a24(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a24_PORTADATAOUT_bus),
	.portbdataout(ram_block3a24_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a24.clk0_core_clock_enable = "ena0";
defparam ram_block3a24.clk1_core_clock_enable = "ena1";
defparam ram_block3a24.data_interleave_offset_in_bits = 1;
defparam ram_block3a24.data_interleave_width_in_bits = 1;
defparam ram_block3a24.init_file = "meminit.hex";
defparam ram_block3a24.init_file_layout = "port_a";
defparam ram_block3a24.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a24.operation_mode = "bidir_dual_port";
defparam ram_block3a24.port_a_address_clear = "none";
defparam ram_block3a24.port_a_address_width = 13;
defparam ram_block3a24.port_a_byte_enable_clock = "none";
defparam ram_block3a24.port_a_data_out_clear = "none";
defparam ram_block3a24.port_a_data_out_clock = "none";
defparam ram_block3a24.port_a_data_width = 1;
defparam ram_block3a24.port_a_first_address = 0;
defparam ram_block3a24.port_a_first_bit_number = 24;
defparam ram_block3a24.port_a_last_address = 8191;
defparam ram_block3a24.port_a_logical_ram_depth = 16384;
defparam ram_block3a24.port_a_logical_ram_width = 32;
defparam ram_block3a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_address_clear = "none";
defparam ram_block3a24.port_b_address_clock = "clock1";
defparam ram_block3a24.port_b_address_width = 13;
defparam ram_block3a24.port_b_data_in_clock = "clock1";
defparam ram_block3a24.port_b_data_out_clear = "none";
defparam ram_block3a24.port_b_data_out_clock = "none";
defparam ram_block3a24.port_b_data_width = 1;
defparam ram_block3a24.port_b_first_address = 0;
defparam ram_block3a24.port_b_first_bit_number = 24;
defparam ram_block3a24.port_b_last_address = 8191;
defparam ram_block3a24.port_b_logical_ram_depth = 16384;
defparam ram_block3a24.port_b_logical_ram_width = 32;
defparam ram_block3a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_read_enable_clock = "clock1";
defparam ram_block3a24.port_b_write_enable_clock = "clock1";
defparam ram_block3a24.ram_block_type = "M9K";
defparam ram_block3a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021830C680DB793600400;
// synopsys translate_on

// Location: M9K_X51_Y33_N0
cycloneive_ram_block ram_block3a57(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a57_PORTADATAOUT_bus),
	.portbdataout(ram_block3a57_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a57.clk0_core_clock_enable = "ena0";
defparam ram_block3a57.clk1_core_clock_enable = "ena1";
defparam ram_block3a57.data_interleave_offset_in_bits = 1;
defparam ram_block3a57.data_interleave_width_in_bits = 1;
defparam ram_block3a57.init_file = "meminit.hex";
defparam ram_block3a57.init_file_layout = "port_a";
defparam ram_block3a57.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a57.operation_mode = "bidir_dual_port";
defparam ram_block3a57.port_a_address_clear = "none";
defparam ram_block3a57.port_a_address_width = 13;
defparam ram_block3a57.port_a_byte_enable_clock = "none";
defparam ram_block3a57.port_a_data_out_clear = "none";
defparam ram_block3a57.port_a_data_out_clock = "none";
defparam ram_block3a57.port_a_data_width = 1;
defparam ram_block3a57.port_a_first_address = 0;
defparam ram_block3a57.port_a_first_bit_number = 25;
defparam ram_block3a57.port_a_last_address = 8191;
defparam ram_block3a57.port_a_logical_ram_depth = 16384;
defparam ram_block3a57.port_a_logical_ram_width = 32;
defparam ram_block3a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_address_clear = "none";
defparam ram_block3a57.port_b_address_clock = "clock1";
defparam ram_block3a57.port_b_address_width = 13;
defparam ram_block3a57.port_b_data_in_clock = "clock1";
defparam ram_block3a57.port_b_data_out_clear = "none";
defparam ram_block3a57.port_b_data_out_clock = "none";
defparam ram_block3a57.port_b_data_width = 1;
defparam ram_block3a57.port_b_first_address = 0;
defparam ram_block3a57.port_b_first_bit_number = 25;
defparam ram_block3a57.port_b_last_address = 8191;
defparam ram_block3a57.port_b_logical_ram_depth = 16384;
defparam ram_block3a57.port_b_logical_ram_width = 32;
defparam ram_block3a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_read_enable_clock = "clock1";
defparam ram_block3a57.port_b_write_enable_clock = "clock1";
defparam ram_block3a57.ram_block_type = "M9K";
defparam ram_block3a57.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y33_N0
cycloneive_ram_block ram_block3a25(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a25_PORTADATAOUT_bus),
	.portbdataout(ram_block3a25_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a25.clk0_core_clock_enable = "ena0";
defparam ram_block3a25.clk1_core_clock_enable = "ena1";
defparam ram_block3a25.data_interleave_offset_in_bits = 1;
defparam ram_block3a25.data_interleave_width_in_bits = 1;
defparam ram_block3a25.init_file = "meminit.hex";
defparam ram_block3a25.init_file_layout = "port_a";
defparam ram_block3a25.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a25.operation_mode = "bidir_dual_port";
defparam ram_block3a25.port_a_address_clear = "none";
defparam ram_block3a25.port_a_address_width = 13;
defparam ram_block3a25.port_a_byte_enable_clock = "none";
defparam ram_block3a25.port_a_data_out_clear = "none";
defparam ram_block3a25.port_a_data_out_clock = "none";
defparam ram_block3a25.port_a_data_width = 1;
defparam ram_block3a25.port_a_first_address = 0;
defparam ram_block3a25.port_a_first_bit_number = 25;
defparam ram_block3a25.port_a_last_address = 8191;
defparam ram_block3a25.port_a_logical_ram_depth = 16384;
defparam ram_block3a25.port_a_logical_ram_width = 32;
defparam ram_block3a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_address_clear = "none";
defparam ram_block3a25.port_b_address_clock = "clock1";
defparam ram_block3a25.port_b_address_width = 13;
defparam ram_block3a25.port_b_data_in_clock = "clock1";
defparam ram_block3a25.port_b_data_out_clear = "none";
defparam ram_block3a25.port_b_data_out_clock = "none";
defparam ram_block3a25.port_b_data_width = 1;
defparam ram_block3a25.port_b_first_address = 0;
defparam ram_block3a25.port_b_first_bit_number = 25;
defparam ram_block3a25.port_b_last_address = 8191;
defparam ram_block3a25.port_b_logical_ram_depth = 16384;
defparam ram_block3a25.port_b_logical_ram_width = 32;
defparam ram_block3a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_read_enable_clock = "clock1";
defparam ram_block3a25.port_b_write_enable_clock = "clock1";
defparam ram_block3a25.ram_block_type = "M9K";
defparam ram_block3a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000CB783600310;
// synopsys translate_on

// Location: M9K_X37_Y29_N0
cycloneive_ram_block ram_block3a58(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a58_PORTADATAOUT_bus),
	.portbdataout(ram_block3a58_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a58.clk0_core_clock_enable = "ena0";
defparam ram_block3a58.clk1_core_clock_enable = "ena1";
defparam ram_block3a58.data_interleave_offset_in_bits = 1;
defparam ram_block3a58.data_interleave_width_in_bits = 1;
defparam ram_block3a58.init_file = "meminit.hex";
defparam ram_block3a58.init_file_layout = "port_a";
defparam ram_block3a58.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a58.operation_mode = "bidir_dual_port";
defparam ram_block3a58.port_a_address_clear = "none";
defparam ram_block3a58.port_a_address_width = 13;
defparam ram_block3a58.port_a_byte_enable_clock = "none";
defparam ram_block3a58.port_a_data_out_clear = "none";
defparam ram_block3a58.port_a_data_out_clock = "none";
defparam ram_block3a58.port_a_data_width = 1;
defparam ram_block3a58.port_a_first_address = 0;
defparam ram_block3a58.port_a_first_bit_number = 26;
defparam ram_block3a58.port_a_last_address = 8191;
defparam ram_block3a58.port_a_logical_ram_depth = 16384;
defparam ram_block3a58.port_a_logical_ram_width = 32;
defparam ram_block3a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_address_clear = "none";
defparam ram_block3a58.port_b_address_clock = "clock1";
defparam ram_block3a58.port_b_address_width = 13;
defparam ram_block3a58.port_b_data_in_clock = "clock1";
defparam ram_block3a58.port_b_data_out_clear = "none";
defparam ram_block3a58.port_b_data_out_clock = "none";
defparam ram_block3a58.port_b_data_width = 1;
defparam ram_block3a58.port_b_first_address = 0;
defparam ram_block3a58.port_b_first_bit_number = 26;
defparam ram_block3a58.port_b_last_address = 8191;
defparam ram_block3a58.port_b_logical_ram_depth = 16384;
defparam ram_block3a58.port_b_logical_ram_width = 32;
defparam ram_block3a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_read_enable_clock = "clock1";
defparam ram_block3a58.port_b_write_enable_clock = "clock1";
defparam ram_block3a58.ram_block_type = "M9K";
defparam ram_block3a58.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y28_N0
cycloneive_ram_block ram_block3a26(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a26_PORTADATAOUT_bus),
	.portbdataout(ram_block3a26_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a26.clk0_core_clock_enable = "ena0";
defparam ram_block3a26.clk1_core_clock_enable = "ena1";
defparam ram_block3a26.data_interleave_offset_in_bits = 1;
defparam ram_block3a26.data_interleave_width_in_bits = 1;
defparam ram_block3a26.init_file = "meminit.hex";
defparam ram_block3a26.init_file_layout = "port_a";
defparam ram_block3a26.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a26.operation_mode = "bidir_dual_port";
defparam ram_block3a26.port_a_address_clear = "none";
defparam ram_block3a26.port_a_address_width = 13;
defparam ram_block3a26.port_a_byte_enable_clock = "none";
defparam ram_block3a26.port_a_data_out_clear = "none";
defparam ram_block3a26.port_a_data_out_clock = "none";
defparam ram_block3a26.port_a_data_width = 1;
defparam ram_block3a26.port_a_first_address = 0;
defparam ram_block3a26.port_a_first_bit_number = 26;
defparam ram_block3a26.port_a_last_address = 8191;
defparam ram_block3a26.port_a_logical_ram_depth = 16384;
defparam ram_block3a26.port_a_logical_ram_width = 32;
defparam ram_block3a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_address_clear = "none";
defparam ram_block3a26.port_b_address_clock = "clock1";
defparam ram_block3a26.port_b_address_width = 13;
defparam ram_block3a26.port_b_data_in_clock = "clock1";
defparam ram_block3a26.port_b_data_out_clear = "none";
defparam ram_block3a26.port_b_data_out_clock = "none";
defparam ram_block3a26.port_b_data_width = 1;
defparam ram_block3a26.port_b_first_address = 0;
defparam ram_block3a26.port_b_first_bit_number = 26;
defparam ram_block3a26.port_b_last_address = 8191;
defparam ram_block3a26.port_b_logical_ram_depth = 16384;
defparam ram_block3a26.port_b_logical_ram_width = 32;
defparam ram_block3a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_read_enable_clock = "clock1";
defparam ram_block3a26.port_b_write_enable_clock = "clock1";
defparam ram_block3a26.ram_block_type = "M9K";
defparam ram_block3a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007CFBDE639B287F0888F;
// synopsys translate_on

// Location: M9K_X37_Y39_N0
cycloneive_ram_block ram_block3a59(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a59_PORTADATAOUT_bus),
	.portbdataout(ram_block3a59_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a59.clk0_core_clock_enable = "ena0";
defparam ram_block3a59.clk1_core_clock_enable = "ena1";
defparam ram_block3a59.data_interleave_offset_in_bits = 1;
defparam ram_block3a59.data_interleave_width_in_bits = 1;
defparam ram_block3a59.init_file = "meminit.hex";
defparam ram_block3a59.init_file_layout = "port_a";
defparam ram_block3a59.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a59.operation_mode = "bidir_dual_port";
defparam ram_block3a59.port_a_address_clear = "none";
defparam ram_block3a59.port_a_address_width = 13;
defparam ram_block3a59.port_a_byte_enable_clock = "none";
defparam ram_block3a59.port_a_data_out_clear = "none";
defparam ram_block3a59.port_a_data_out_clock = "none";
defparam ram_block3a59.port_a_data_width = 1;
defparam ram_block3a59.port_a_first_address = 0;
defparam ram_block3a59.port_a_first_bit_number = 27;
defparam ram_block3a59.port_a_last_address = 8191;
defparam ram_block3a59.port_a_logical_ram_depth = 16384;
defparam ram_block3a59.port_a_logical_ram_width = 32;
defparam ram_block3a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_address_clear = "none";
defparam ram_block3a59.port_b_address_clock = "clock1";
defparam ram_block3a59.port_b_address_width = 13;
defparam ram_block3a59.port_b_data_in_clock = "clock1";
defparam ram_block3a59.port_b_data_out_clear = "none";
defparam ram_block3a59.port_b_data_out_clock = "none";
defparam ram_block3a59.port_b_data_width = 1;
defparam ram_block3a59.port_b_first_address = 0;
defparam ram_block3a59.port_b_first_bit_number = 27;
defparam ram_block3a59.port_b_last_address = 8191;
defparam ram_block3a59.port_b_logical_ram_depth = 16384;
defparam ram_block3a59.port_b_logical_ram_width = 32;
defparam ram_block3a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_read_enable_clock = "clock1";
defparam ram_block3a59.port_b_write_enable_clock = "clock1";
defparam ram_block3a59.ram_block_type = "M9K";
defparam ram_block3a59.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y37_N0
cycloneive_ram_block ram_block3a27(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a27_PORTADATAOUT_bus),
	.portbdataout(ram_block3a27_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a27.clk0_core_clock_enable = "ena0";
defparam ram_block3a27.clk1_core_clock_enable = "ena1";
defparam ram_block3a27.data_interleave_offset_in_bits = 1;
defparam ram_block3a27.data_interleave_width_in_bits = 1;
defparam ram_block3a27.init_file = "meminit.hex";
defparam ram_block3a27.init_file_layout = "port_a";
defparam ram_block3a27.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a27.operation_mode = "bidir_dual_port";
defparam ram_block3a27.port_a_address_clear = "none";
defparam ram_block3a27.port_a_address_width = 13;
defparam ram_block3a27.port_a_byte_enable_clock = "none";
defparam ram_block3a27.port_a_data_out_clear = "none";
defparam ram_block3a27.port_a_data_out_clock = "none";
defparam ram_block3a27.port_a_data_width = 1;
defparam ram_block3a27.port_a_first_address = 0;
defparam ram_block3a27.port_a_first_bit_number = 27;
defparam ram_block3a27.port_a_last_address = 8191;
defparam ram_block3a27.port_a_logical_ram_depth = 16384;
defparam ram_block3a27.port_a_logical_ram_width = 32;
defparam ram_block3a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_address_clear = "none";
defparam ram_block3a27.port_b_address_clock = "clock1";
defparam ram_block3a27.port_b_address_width = 13;
defparam ram_block3a27.port_b_data_in_clock = "clock1";
defparam ram_block3a27.port_b_data_out_clear = "none";
defparam ram_block3a27.port_b_data_out_clock = "none";
defparam ram_block3a27.port_b_data_width = 1;
defparam ram_block3a27.port_b_first_address = 0;
defparam ram_block3a27.port_b_first_bit_number = 27;
defparam ram_block3a27.port_b_last_address = 8191;
defparam ram_block3a27.port_b_logical_ram_depth = 16384;
defparam ram_block3a27.port_b_logical_ram_width = 32;
defparam ram_block3a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_read_enable_clock = "clock1";
defparam ram_block3a27.port_b_write_enable_clock = "clock1";
defparam ram_block3a27.ram_block_type = "M9K";
defparam ram_block3a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010E1C6264AD282C08088;
// synopsys translate_on

// Location: M9K_X37_Y32_N0
cycloneive_ram_block ram_block3a60(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a60_PORTADATAOUT_bus),
	.portbdataout(ram_block3a60_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a60.clk0_core_clock_enable = "ena0";
defparam ram_block3a60.clk1_core_clock_enable = "ena1";
defparam ram_block3a60.data_interleave_offset_in_bits = 1;
defparam ram_block3a60.data_interleave_width_in_bits = 1;
defparam ram_block3a60.init_file = "meminit.hex";
defparam ram_block3a60.init_file_layout = "port_a";
defparam ram_block3a60.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a60.operation_mode = "bidir_dual_port";
defparam ram_block3a60.port_a_address_clear = "none";
defparam ram_block3a60.port_a_address_width = 13;
defparam ram_block3a60.port_a_byte_enable_clock = "none";
defparam ram_block3a60.port_a_data_out_clear = "none";
defparam ram_block3a60.port_a_data_out_clock = "none";
defparam ram_block3a60.port_a_data_width = 1;
defparam ram_block3a60.port_a_first_address = 0;
defparam ram_block3a60.port_a_first_bit_number = 28;
defparam ram_block3a60.port_a_last_address = 8191;
defparam ram_block3a60.port_a_logical_ram_depth = 16384;
defparam ram_block3a60.port_a_logical_ram_width = 32;
defparam ram_block3a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_address_clear = "none";
defparam ram_block3a60.port_b_address_clock = "clock1";
defparam ram_block3a60.port_b_address_width = 13;
defparam ram_block3a60.port_b_data_in_clock = "clock1";
defparam ram_block3a60.port_b_data_out_clear = "none";
defparam ram_block3a60.port_b_data_out_clock = "none";
defparam ram_block3a60.port_b_data_width = 1;
defparam ram_block3a60.port_b_first_address = 0;
defparam ram_block3a60.port_b_first_bit_number = 28;
defparam ram_block3a60.port_b_last_address = 8191;
defparam ram_block3a60.port_b_logical_ram_depth = 16384;
defparam ram_block3a60.port_b_logical_ram_width = 32;
defparam ram_block3a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_read_enable_clock = "clock1";
defparam ram_block3a60.port_b_write_enable_clock = "clock1";
defparam ram_block3a60.ram_block_type = "M9K";
defparam ram_block3a60.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y30_N0
cycloneive_ram_block ram_block3a28(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a28_PORTADATAOUT_bus),
	.portbdataout(ram_block3a28_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a28.clk0_core_clock_enable = "ena0";
defparam ram_block3a28.clk1_core_clock_enable = "ena1";
defparam ram_block3a28.data_interleave_offset_in_bits = 1;
defparam ram_block3a28.data_interleave_width_in_bits = 1;
defparam ram_block3a28.init_file = "meminit.hex";
defparam ram_block3a28.init_file_layout = "port_a";
defparam ram_block3a28.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a28.operation_mode = "bidir_dual_port";
defparam ram_block3a28.port_a_address_clear = "none";
defparam ram_block3a28.port_a_address_width = 13;
defparam ram_block3a28.port_a_byte_enable_clock = "none";
defparam ram_block3a28.port_a_data_out_clear = "none";
defparam ram_block3a28.port_a_data_out_clock = "none";
defparam ram_block3a28.port_a_data_width = 1;
defparam ram_block3a28.port_a_first_address = 0;
defparam ram_block3a28.port_a_first_bit_number = 28;
defparam ram_block3a28.port_a_last_address = 8191;
defparam ram_block3a28.port_a_logical_ram_depth = 16384;
defparam ram_block3a28.port_a_logical_ram_width = 32;
defparam ram_block3a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_address_clear = "none";
defparam ram_block3a28.port_b_address_clock = "clock1";
defparam ram_block3a28.port_b_address_width = 13;
defparam ram_block3a28.port_b_data_in_clock = "clock1";
defparam ram_block3a28.port_b_data_out_clear = "none";
defparam ram_block3a28.port_b_data_out_clock = "none";
defparam ram_block3a28.port_b_data_width = 1;
defparam ram_block3a28.port_b_first_address = 0;
defparam ram_block3a28.port_b_first_bit_number = 28;
defparam ram_block3a28.port_b_last_address = 8191;
defparam ram_block3a28.port_b_logical_ram_depth = 16384;
defparam ram_block3a28.port_b_logical_ram_width = 32;
defparam ram_block3a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_read_enable_clock = "clock1";
defparam ram_block3a28.port_b_write_enable_clock = "clock1";
defparam ram_block3a28.ram_block_type = "M9K";
defparam ram_block3a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008100011B00926100807;
// synopsys translate_on

// Location: M9K_X64_Y28_N0
cycloneive_ram_block ram_block3a61(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a61_PORTADATAOUT_bus),
	.portbdataout(ram_block3a61_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a61.clk0_core_clock_enable = "ena0";
defparam ram_block3a61.clk1_core_clock_enable = "ena1";
defparam ram_block3a61.data_interleave_offset_in_bits = 1;
defparam ram_block3a61.data_interleave_width_in_bits = 1;
defparam ram_block3a61.init_file = "meminit.hex";
defparam ram_block3a61.init_file_layout = "port_a";
defparam ram_block3a61.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a61.operation_mode = "bidir_dual_port";
defparam ram_block3a61.port_a_address_clear = "none";
defparam ram_block3a61.port_a_address_width = 13;
defparam ram_block3a61.port_a_byte_enable_clock = "none";
defparam ram_block3a61.port_a_data_out_clear = "none";
defparam ram_block3a61.port_a_data_out_clock = "none";
defparam ram_block3a61.port_a_data_width = 1;
defparam ram_block3a61.port_a_first_address = 0;
defparam ram_block3a61.port_a_first_bit_number = 29;
defparam ram_block3a61.port_a_last_address = 8191;
defparam ram_block3a61.port_a_logical_ram_depth = 16384;
defparam ram_block3a61.port_a_logical_ram_width = 32;
defparam ram_block3a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_address_clear = "none";
defparam ram_block3a61.port_b_address_clock = "clock1";
defparam ram_block3a61.port_b_address_width = 13;
defparam ram_block3a61.port_b_data_in_clock = "clock1";
defparam ram_block3a61.port_b_data_out_clear = "none";
defparam ram_block3a61.port_b_data_out_clock = "none";
defparam ram_block3a61.port_b_data_width = 1;
defparam ram_block3a61.port_b_first_address = 0;
defparam ram_block3a61.port_b_first_bit_number = 29;
defparam ram_block3a61.port_b_last_address = 8191;
defparam ram_block3a61.port_b_logical_ram_depth = 16384;
defparam ram_block3a61.port_b_logical_ram_width = 32;
defparam ram_block3a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_read_enable_clock = "clock1";
defparam ram_block3a61.port_b_write_enable_clock = "clock1";
defparam ram_block3a61.ram_block_type = "M9K";
defparam ram_block3a61.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y25_N0
cycloneive_ram_block ram_block3a29(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a29_PORTADATAOUT_bus),
	.portbdataout(ram_block3a29_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a29.clk0_core_clock_enable = "ena0";
defparam ram_block3a29.clk1_core_clock_enable = "ena1";
defparam ram_block3a29.data_interleave_offset_in_bits = 1;
defparam ram_block3a29.data_interleave_width_in_bits = 1;
defparam ram_block3a29.init_file = "meminit.hex";
defparam ram_block3a29.init_file_layout = "port_a";
defparam ram_block3a29.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a29.operation_mode = "bidir_dual_port";
defparam ram_block3a29.port_a_address_clear = "none";
defparam ram_block3a29.port_a_address_width = 13;
defparam ram_block3a29.port_a_byte_enable_clock = "none";
defparam ram_block3a29.port_a_data_out_clear = "none";
defparam ram_block3a29.port_a_data_out_clock = "none";
defparam ram_block3a29.port_a_data_width = 1;
defparam ram_block3a29.port_a_first_address = 0;
defparam ram_block3a29.port_a_first_bit_number = 29;
defparam ram_block3a29.port_a_last_address = 8191;
defparam ram_block3a29.port_a_logical_ram_depth = 16384;
defparam ram_block3a29.port_a_logical_ram_width = 32;
defparam ram_block3a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_address_clear = "none";
defparam ram_block3a29.port_b_address_clock = "clock1";
defparam ram_block3a29.port_b_address_width = 13;
defparam ram_block3a29.port_b_data_in_clock = "clock1";
defparam ram_block3a29.port_b_data_out_clear = "none";
defparam ram_block3a29.port_b_data_out_clock = "none";
defparam ram_block3a29.port_b_data_width = 1;
defparam ram_block3a29.port_b_first_address = 0;
defparam ram_block3a29.port_b_first_bit_number = 29;
defparam ram_block3a29.port_b_last_address = 8191;
defparam ram_block3a29.port_b_logical_ram_depth = 16384;
defparam ram_block3a29.port_b_logical_ram_width = 32;
defparam ram_block3a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_read_enable_clock = "clock1";
defparam ram_block3a29.port_b_write_enable_clock = "clock1";
defparam ram_block3a29.ram_block_type = "M9K";
defparam ram_block3a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000078F3DE001B007700807;
// synopsys translate_on

// Location: M9K_X78_Y29_N0
cycloneive_ram_block ram_block3a62(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a62_PORTADATAOUT_bus),
	.portbdataout(ram_block3a62_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a62.clk0_core_clock_enable = "ena0";
defparam ram_block3a62.clk1_core_clock_enable = "ena1";
defparam ram_block3a62.data_interleave_offset_in_bits = 1;
defparam ram_block3a62.data_interleave_width_in_bits = 1;
defparam ram_block3a62.init_file = "meminit.hex";
defparam ram_block3a62.init_file_layout = "port_a";
defparam ram_block3a62.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a62.operation_mode = "bidir_dual_port";
defparam ram_block3a62.port_a_address_clear = "none";
defparam ram_block3a62.port_a_address_width = 13;
defparam ram_block3a62.port_a_byte_enable_clock = "none";
defparam ram_block3a62.port_a_data_out_clear = "none";
defparam ram_block3a62.port_a_data_out_clock = "none";
defparam ram_block3a62.port_a_data_width = 1;
defparam ram_block3a62.port_a_first_address = 0;
defparam ram_block3a62.port_a_first_bit_number = 30;
defparam ram_block3a62.port_a_last_address = 8191;
defparam ram_block3a62.port_a_logical_ram_depth = 16384;
defparam ram_block3a62.port_a_logical_ram_width = 32;
defparam ram_block3a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_address_clear = "none";
defparam ram_block3a62.port_b_address_clock = "clock1";
defparam ram_block3a62.port_b_address_width = 13;
defparam ram_block3a62.port_b_data_in_clock = "clock1";
defparam ram_block3a62.port_b_data_out_clear = "none";
defparam ram_block3a62.port_b_data_out_clock = "none";
defparam ram_block3a62.port_b_data_width = 1;
defparam ram_block3a62.port_b_first_address = 0;
defparam ram_block3a62.port_b_first_bit_number = 30;
defparam ram_block3a62.port_b_last_address = 8191;
defparam ram_block3a62.port_b_logical_ram_depth = 16384;
defparam ram_block3a62.port_b_logical_ram_width = 32;
defparam ram_block3a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_read_enable_clock = "clock1";
defparam ram_block3a62.port_b_write_enable_clock = "clock1";
defparam ram_block3a62.ram_block_type = "M9K";
defparam ram_block3a62.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y28_N0
cycloneive_ram_block ram_block3a30(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a30_PORTADATAOUT_bus),
	.portbdataout(ram_block3a30_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a30.clk0_core_clock_enable = "ena0";
defparam ram_block3a30.clk1_core_clock_enable = "ena1";
defparam ram_block3a30.data_interleave_offset_in_bits = 1;
defparam ram_block3a30.data_interleave_width_in_bits = 1;
defparam ram_block3a30.init_file = "meminit.hex";
defparam ram_block3a30.init_file_layout = "port_a";
defparam ram_block3a30.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a30.operation_mode = "bidir_dual_port";
defparam ram_block3a30.port_a_address_clear = "none";
defparam ram_block3a30.port_a_address_width = 13;
defparam ram_block3a30.port_a_byte_enable_clock = "none";
defparam ram_block3a30.port_a_data_out_clear = "none";
defparam ram_block3a30.port_a_data_out_clock = "none";
defparam ram_block3a30.port_a_data_width = 1;
defparam ram_block3a30.port_a_first_address = 0;
defparam ram_block3a30.port_a_first_bit_number = 30;
defparam ram_block3a30.port_a_last_address = 8191;
defparam ram_block3a30.port_a_logical_ram_depth = 16384;
defparam ram_block3a30.port_a_logical_ram_width = 32;
defparam ram_block3a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_address_clear = "none";
defparam ram_block3a30.port_b_address_clock = "clock1";
defparam ram_block3a30.port_b_address_width = 13;
defparam ram_block3a30.port_b_data_in_clock = "clock1";
defparam ram_block3a30.port_b_data_out_clear = "none";
defparam ram_block3a30.port_b_data_out_clock = "none";
defparam ram_block3a30.port_b_data_width = 1;
defparam ram_block3a30.port_b_first_address = 0;
defparam ram_block3a30.port_b_first_bit_number = 30;
defparam ram_block3a30.port_b_last_address = 8191;
defparam ram_block3a30.port_b_logical_ram_depth = 16384;
defparam ram_block3a30.port_b_logical_ram_width = 32;
defparam ram_block3a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_read_enable_clock = "clock1";
defparam ram_block3a30.port_b_write_enable_clock = "clock1";
defparam ram_block3a30.ram_block_type = "M9K";
defparam ram_block3a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000;
// synopsys translate_on

// Location: M9K_X78_Y32_N0
cycloneive_ram_block ram_block3a63(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a63_PORTADATAOUT_bus),
	.portbdataout(ram_block3a63_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a63.clk0_core_clock_enable = "ena0";
defparam ram_block3a63.clk1_core_clock_enable = "ena1";
defparam ram_block3a63.data_interleave_offset_in_bits = 1;
defparam ram_block3a63.data_interleave_width_in_bits = 1;
defparam ram_block3a63.init_file = "meminit.hex";
defparam ram_block3a63.init_file_layout = "port_a";
defparam ram_block3a63.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a63.operation_mode = "bidir_dual_port";
defparam ram_block3a63.port_a_address_clear = "none";
defparam ram_block3a63.port_a_address_width = 13;
defparam ram_block3a63.port_a_byte_enable_clock = "none";
defparam ram_block3a63.port_a_data_out_clear = "none";
defparam ram_block3a63.port_a_data_out_clock = "none";
defparam ram_block3a63.port_a_data_width = 1;
defparam ram_block3a63.port_a_first_address = 0;
defparam ram_block3a63.port_a_first_bit_number = 31;
defparam ram_block3a63.port_a_last_address = 8191;
defparam ram_block3a63.port_a_logical_ram_depth = 16384;
defparam ram_block3a63.port_a_logical_ram_width = 32;
defparam ram_block3a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_address_clear = "none";
defparam ram_block3a63.port_b_address_clock = "clock1";
defparam ram_block3a63.port_b_address_width = 13;
defparam ram_block3a63.port_b_data_in_clock = "clock1";
defparam ram_block3a63.port_b_data_out_clear = "none";
defparam ram_block3a63.port_b_data_out_clock = "none";
defparam ram_block3a63.port_b_data_width = 1;
defparam ram_block3a63.port_b_first_address = 0;
defparam ram_block3a63.port_b_first_bit_number = 31;
defparam ram_block3a63.port_b_last_address = 8191;
defparam ram_block3a63.port_b_logical_ram_depth = 16384;
defparam ram_block3a63.port_b_logical_ram_width = 32;
defparam ram_block3a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_read_enable_clock = "clock1";
defparam ram_block3a63.port_b_write_enable_clock = "clock1";
defparam ram_block3a63.ram_block_type = "M9K";
defparam ram_block3a63.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y34_N0
cycloneive_ram_block ram_block3a31(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a31_PORTADATAOUT_bus),
	.portbdataout(ram_block3a31_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a31.clk0_core_clock_enable = "ena0";
defparam ram_block3a31.clk1_core_clock_enable = "ena1";
defparam ram_block3a31.data_interleave_offset_in_bits = 1;
defparam ram_block3a31.data_interleave_width_in_bits = 1;
defparam ram_block3a31.init_file = "meminit.hex";
defparam ram_block3a31.init_file_layout = "port_a";
defparam ram_block3a31.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a31.operation_mode = "bidir_dual_port";
defparam ram_block3a31.port_a_address_clear = "none";
defparam ram_block3a31.port_a_address_width = 13;
defparam ram_block3a31.port_a_byte_enable_clock = "none";
defparam ram_block3a31.port_a_data_out_clear = "none";
defparam ram_block3a31.port_a_data_out_clock = "none";
defparam ram_block3a31.port_a_data_width = 1;
defparam ram_block3a31.port_a_first_address = 0;
defparam ram_block3a31.port_a_first_bit_number = 31;
defparam ram_block3a31.port_a_last_address = 8191;
defparam ram_block3a31.port_a_logical_ram_depth = 16384;
defparam ram_block3a31.port_a_logical_ram_width = 32;
defparam ram_block3a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_address_clear = "none";
defparam ram_block3a31.port_b_address_clock = "clock1";
defparam ram_block3a31.port_b_address_width = 13;
defparam ram_block3a31.port_b_data_in_clock = "clock1";
defparam ram_block3a31.port_b_data_out_clear = "none";
defparam ram_block3a31.port_b_data_out_clock = "none";
defparam ram_block3a31.port_b_data_width = 1;
defparam ram_block3a31.port_b_first_address = 0;
defparam ram_block3a31.port_b_first_bit_number = 31;
defparam ram_block3a31.port_b_last_address = 8191;
defparam ram_block3a31.port_b_logical_ram_depth = 16384;
defparam ram_block3a31.port_b_logical_ram_width = 32;
defparam ram_block3a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_read_enable_clock = "clock1";
defparam ram_block3a31.port_b_write_enable_clock = "clock1";
defparam ram_block3a31.ram_block_type = "M9K";
defparam ram_block3a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000C18426089282400008;
// synopsys translate_on

// Location: FF_X57_Y38_N29
dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_a_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N21
dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(\address_reg_b[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_b_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N20
cycloneive_lcell_comb \address_reg_b[0]~feeder (
// Equation(s):
// \address_reg_b[0]~feeder_combout  = ram_rom_addr_reg_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_13),
	.cin(gnd),
	.combout(\address_reg_b[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \address_reg_b[0]~feeder .lut_mask = 16'hFF00;
defparam \address_reg_b[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa (
	ramaddr,
	ramWEN,
	always1,
	eq_node_1,
	eq_node_0,
	devpor,
	devclrn,
	devoe);
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	eq_node_1;
output 	eq_node_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X61_Y38_N30
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (!\ramWEN~0_combout  & (!\ramaddr~29_combout  & always1))

	.dataa(ramWEN),
	.datab(gnd),
	.datac(ramaddr),
	.datad(always1),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h0500;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N0
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (!\ramWEN~0_combout  & (\ramaddr~29_combout  & always1))

	.dataa(ramWEN),
	.datab(gnd),
	.datac(ramaddr),
	.datad(always1),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h5000;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa_1 (
	ram_rom_addr_reg_13,
	sdr,
	eq_node_1,
	eq_node_0,
	irf_reg_2_1,
	state_5,
	devpor,
	devclrn,
	devoe);
input 	ram_rom_addr_reg_13;
input 	sdr;
output 	eq_node_1;
output 	eq_node_0;
input 	irf_reg_2_1;
input 	state_5;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X46_Y34_N16
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & (sdr & (ram_rom_addr_reg_13 & \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q )))

	.dataa(state_5),
	.datab(sdr),
	.datac(ram_rom_addr_reg_13),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h8000;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N10
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & (sdr & (!ram_rom_addr_reg_13 & \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q )))

	.dataa(state_5),
	.datab(sdr),
	.datac(ram_rom_addr_reg_13),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h0800;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_mod_ram_rom (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg1,
	ram_rom_data_reg_0,
	ram_rom_addr_reg_13,
	ram_rom_addr_reg_0,
	ram_rom_addr_reg_1,
	ram_rom_addr_reg_2,
	ram_rom_addr_reg_3,
	ram_rom_addr_reg_4,
	ram_rom_addr_reg_5,
	ram_rom_addr_reg_6,
	ram_rom_addr_reg_7,
	ram_rom_addr_reg_8,
	ram_rom_addr_reg_9,
	ram_rom_addr_reg_10,
	ram_rom_addr_reg_11,
	ram_rom_addr_reg_12,
	ram_rom_data_reg_1,
	ram_rom_data_reg_2,
	ram_rom_data_reg_3,
	ram_rom_data_reg_4,
	ram_rom_data_reg_5,
	ram_rom_data_reg_6,
	ram_rom_data_reg_7,
	ram_rom_data_reg_8,
	ram_rom_data_reg_9,
	ram_rom_data_reg_10,
	ram_rom_data_reg_11,
	ram_rom_data_reg_12,
	ram_rom_data_reg_13,
	ram_rom_data_reg_14,
	ram_rom_data_reg_15,
	ram_rom_data_reg_16,
	ram_rom_data_reg_17,
	ram_rom_data_reg_18,
	ram_rom_data_reg_19,
	ram_rom_data_reg_20,
	ram_rom_data_reg_21,
	ram_rom_data_reg_22,
	ram_rom_data_reg_23,
	ram_rom_data_reg_24,
	ram_rom_data_reg_25,
	ram_rom_data_reg_26,
	ram_rom_data_reg_27,
	ram_rom_data_reg_28,
	ram_rom_data_reg_29,
	ram_rom_data_reg_30,
	ram_rom_data_reg_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	sdr,
	address_reg_b_0,
	altera_internal_jtag,
	state_4,
	ir_in,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_4_1,
	node_ena_1,
	clr,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	raw_tck,
	devpor,
	devclrn,
	devoe);
input 	ram_block3a32;
input 	ram_block3a0;
input 	ram_block3a33;
input 	ram_block3a1;
input 	ram_block3a34;
input 	ram_block3a2;
input 	ram_block3a35;
input 	ram_block3a3;
input 	ram_block3a36;
input 	ram_block3a4;
input 	ram_block3a37;
input 	ram_block3a5;
input 	ram_block3a38;
input 	ram_block3a6;
input 	ram_block3a39;
input 	ram_block3a7;
input 	ram_block3a40;
input 	ram_block3a8;
input 	ram_block3a41;
input 	ram_block3a9;
input 	ram_block3a42;
input 	ram_block3a10;
input 	ram_block3a43;
input 	ram_block3a11;
input 	ram_block3a44;
input 	ram_block3a12;
input 	ram_block3a45;
input 	ram_block3a13;
input 	ram_block3a46;
input 	ram_block3a14;
input 	ram_block3a47;
input 	ram_block3a15;
input 	ram_block3a48;
input 	ram_block3a16;
input 	ram_block3a49;
input 	ram_block3a17;
input 	ram_block3a50;
input 	ram_block3a18;
input 	ram_block3a51;
input 	ram_block3a19;
input 	ram_block3a52;
input 	ram_block3a20;
input 	ram_block3a53;
input 	ram_block3a21;
input 	ram_block3a54;
input 	ram_block3a22;
input 	ram_block3a55;
input 	ram_block3a23;
input 	ram_block3a56;
input 	ram_block3a24;
input 	ram_block3a57;
input 	ram_block3a25;
input 	ram_block3a58;
input 	ram_block3a26;
input 	ram_block3a59;
input 	ram_block3a27;
input 	ram_block3a60;
input 	ram_block3a28;
input 	ram_block3a61;
input 	ram_block3a29;
input 	ram_block3a62;
input 	ram_block3a30;
input 	ram_block3a63;
input 	ram_block3a31;
output 	is_in_use_reg1;
output 	ram_rom_data_reg_0;
output 	ram_rom_addr_reg_13;
output 	ram_rom_addr_reg_0;
output 	ram_rom_addr_reg_1;
output 	ram_rom_addr_reg_2;
output 	ram_rom_addr_reg_3;
output 	ram_rom_addr_reg_4;
output 	ram_rom_addr_reg_5;
output 	ram_rom_addr_reg_6;
output 	ram_rom_addr_reg_7;
output 	ram_rom_addr_reg_8;
output 	ram_rom_addr_reg_9;
output 	ram_rom_addr_reg_10;
output 	ram_rom_addr_reg_11;
output 	ram_rom_addr_reg_12;
output 	ram_rom_data_reg_1;
output 	ram_rom_data_reg_2;
output 	ram_rom_data_reg_3;
output 	ram_rom_data_reg_4;
output 	ram_rom_data_reg_5;
output 	ram_rom_data_reg_6;
output 	ram_rom_data_reg_7;
output 	ram_rom_data_reg_8;
output 	ram_rom_data_reg_9;
output 	ram_rom_data_reg_10;
output 	ram_rom_data_reg_11;
output 	ram_rom_data_reg_12;
output 	ram_rom_data_reg_13;
output 	ram_rom_data_reg_14;
output 	ram_rom_data_reg_15;
output 	ram_rom_data_reg_16;
output 	ram_rom_data_reg_17;
output 	ram_rom_data_reg_18;
output 	ram_rom_data_reg_19;
output 	ram_rom_data_reg_20;
output 	ram_rom_data_reg_21;
output 	ram_rom_data_reg_22;
output 	ram_rom_data_reg_23;
output 	ram_rom_data_reg_24;
output 	ram_rom_data_reg_25;
output 	ram_rom_data_reg_26;
output 	ram_rom_data_reg_27;
output 	ram_rom_data_reg_28;
output 	ram_rom_data_reg_29;
output 	ram_rom_data_reg_30;
output 	ram_rom_data_reg_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
output 	sdr;
input 	address_reg_b_0;
input 	altera_internal_jtag;
input 	state_4;
input 	[4:0] ir_in;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	raw_tck;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~6_combout ;
wire \ram_rom_data_shift_cntr_reg[3]~8_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~12_combout ;
wire \is_in_use_reg~0_combout ;
wire \ram_rom_data_reg[0]~0_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \ram_rom_data_shift_cntr_reg[1]~5_combout ;
wire \Add1~3 ;
wire \Add1~4_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~4_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~11_combout ;
wire \ram_rom_data_shift_cntr_reg[2]~9_combout ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~8_combout ;
wire \ram_rom_data_shift_cntr_reg[4]~7_combout ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~10_combout ;
wire \Equal1~0_combout ;
wire \Add1~0_combout ;
wire \ram_rom_data_shift_cntr_reg[0]~6_combout ;
wire \Equal1~1_combout ;
wire \process_0~2_combout ;
wire \ram_rom_data_reg[0]~32_combout ;
wire \ram_rom_addr_reg[0]~15 ;
wire \ram_rom_addr_reg[1]~17 ;
wire \ram_rom_addr_reg[2]~19 ;
wire \ram_rom_addr_reg[3]~21 ;
wire \ram_rom_addr_reg[4]~23 ;
wire \ram_rom_addr_reg[5]~25 ;
wire \ram_rom_addr_reg[6]~27 ;
wire \ram_rom_addr_reg[7]~29 ;
wire \ram_rom_addr_reg[8]~31 ;
wire \ram_rom_addr_reg[9]~33 ;
wire \ram_rom_addr_reg[10]~35 ;
wire \ram_rom_addr_reg[11]~37 ;
wire \ram_rom_addr_reg[12]~39 ;
wire \ram_rom_addr_reg[13]~40_combout ;
wire \process_0~3_combout ;
wire \ram_rom_addr_reg[9]~42_combout ;
wire \ram_rom_addr_reg[9]~43_combout ;
wire \ram_rom_addr_reg[0]~14_combout ;
wire \ram_rom_addr_reg[1]~16_combout ;
wire \ram_rom_addr_reg[2]~18_combout ;
wire \ram_rom_addr_reg[3]~20_combout ;
wire \ram_rom_addr_reg[4]~22_combout ;
wire \ram_rom_addr_reg[5]~24_combout ;
wire \ram_rom_addr_reg[6]~26_combout ;
wire \ram_rom_addr_reg[7]~28_combout ;
wire \ram_rom_addr_reg[8]~30_combout ;
wire \ram_rom_addr_reg[9]~32_combout ;
wire \ram_rom_addr_reg[10]~34_combout ;
wire \ram_rom_addr_reg[11]~36_combout ;
wire \ram_rom_addr_reg[12]~38_combout ;
wire \ram_rom_data_reg[1]~1_combout ;
wire \ram_rom_data_reg[2]~2_combout ;
wire \ram_rom_data_reg[3]~3_combout ;
wire \ram_rom_data_reg[4]~4_combout ;
wire \ram_rom_data_reg[5]~5_combout ;
wire \ram_rom_data_reg[6]~6_combout ;
wire \ram_rom_data_reg[7]~7_combout ;
wire \ram_rom_data_reg[8]~8_combout ;
wire \ram_rom_data_reg[9]~9_combout ;
wire \ram_rom_data_reg[10]~10_combout ;
wire \ram_rom_data_reg[11]~11_combout ;
wire \ram_rom_data_reg[12]~12_combout ;
wire \ram_rom_data_reg[13]~13_combout ;
wire \ram_rom_data_reg[14]~14_combout ;
wire \ram_rom_data_reg[15]~15_combout ;
wire \ram_rom_data_reg[16]~16_combout ;
wire \ram_rom_data_reg[17]~17_combout ;
wire \ram_rom_data_reg[18]~18_combout ;
wire \ram_rom_data_reg[19]~19_combout ;
wire \ram_rom_data_reg[20]~20_combout ;
wire \ram_rom_data_reg[21]~21_combout ;
wire \ram_rom_data_reg[22]~22_combout ;
wire \ram_rom_data_reg[23]~23_combout ;
wire \ram_rom_data_reg[24]~24_combout ;
wire \ram_rom_data_reg[25]~25_combout ;
wire \ram_rom_data_reg[26]~26_combout ;
wire \ram_rom_data_reg[27]~27_combout ;
wire \ram_rom_data_reg[28]~28_combout ;
wire \ram_rom_data_reg[29]~29_combout ;
wire \ram_rom_data_reg[30]~30_combout ;
wire \ram_rom_data_reg[31]~31_combout ;
wire \ir_loaded_address_reg[0]~feeder_combout ;
wire \process_0~0_combout ;
wire \process_0~1_combout ;
wire \ir_loaded_address_reg[1]~feeder_combout ;
wire \ir_loaded_address_reg[2]~feeder_combout ;
wire \ir_loaded_address_reg[3]~feeder_combout ;
wire \bypass_reg_out~0_combout ;
wire \bypass_reg_out~q ;
wire \tdo~0_combout ;
wire [5:0] ram_rom_data_shift_cntr_reg;
wire [3:0] \ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR ;


sld_rom_sr \ram_rom_logic_gen:name_gen:info_rom_sr (
	.WORD_SR_0(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.sdr(sdr),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.TCK(raw_tck),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X47_Y34_N14
cycloneive_lcell_comb \Add1~6 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X47_Y34_N7
dffeas \ram_rom_data_shift_cntr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[3]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N6
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[3]~8 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~6_combout ),
	.datac(ram_rom_data_shift_cntr_reg[3]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3]~8 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N30
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~12 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(\Equal1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~12 .lut_mask = 16'h80FF;
defparam \ram_rom_data_shift_cntr_reg[5]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N13
dffeas is_in_use_reg(
	.clk(raw_tck),
	.d(\is_in_use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(ir_in[0]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(is_in_use_reg1),
	.prn(vcc));
// synopsys translate_off
defparam is_in_use_reg.is_wysiwyg = "true";
defparam is_in_use_reg.power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N1
dffeas \ram_rom_data_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[0]~0_combout ),
	.asdata(ram_rom_data_reg_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N31
dffeas \ram_rom_addr_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[13]~40_combout ),
	.asdata(altera_internal_jtag),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N5
dffeas \ram_rom_addr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[0]~14_combout ),
	.asdata(ram_rom_addr_reg_1),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N7
dffeas \ram_rom_addr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[1]~16_combout ),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N9
dffeas \ram_rom_addr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[2]~18_combout ),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N11
dffeas \ram_rom_addr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[3]~20_combout ),
	.asdata(ram_rom_addr_reg_4),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N13
dffeas \ram_rom_addr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[4]~22_combout ),
	.asdata(ram_rom_addr_reg_5),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N15
dffeas \ram_rom_addr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[5]~24_combout ),
	.asdata(ram_rom_addr_reg_6),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N17
dffeas \ram_rom_addr_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[6]~26_combout ),
	.asdata(ram_rom_addr_reg_7),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N19
dffeas \ram_rom_addr_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[7]~28_combout ),
	.asdata(ram_rom_addr_reg_8),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N21
dffeas \ram_rom_addr_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[8]~30_combout ),
	.asdata(ram_rom_addr_reg_9),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N23
dffeas \ram_rom_addr_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[9]~32_combout ),
	.asdata(ram_rom_addr_reg_10),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N25
dffeas \ram_rom_addr_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[10]~34_combout ),
	.asdata(ram_rom_addr_reg_11),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N27
dffeas \ram_rom_addr_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[11]~36_combout ),
	.asdata(ram_rom_addr_reg_12),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N29
dffeas \ram_rom_addr_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[12]~38_combout ),
	.asdata(ram_rom_addr_reg_13),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[9]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N17
dffeas \ram_rom_data_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[1]~1_combout ),
	.asdata(ram_rom_data_reg_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N23
dffeas \ram_rom_data_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[2]~2_combout ),
	.asdata(ram_rom_data_reg_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N9
dffeas \ram_rom_data_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[3]~3_combout ),
	.asdata(ram_rom_data_reg_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N27
dffeas \ram_rom_data_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[4]~4_combout ),
	.asdata(ram_rom_data_reg_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N25
dffeas \ram_rom_data_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[5]~5_combout ),
	.asdata(ram_rom_data_reg_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N15
dffeas \ram_rom_data_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[6]~6_combout ),
	.asdata(ram_rom_data_reg_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N21
dffeas \ram_rom_data_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[7]~7_combout ),
	.asdata(ram_rom_data_reg_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N31
dffeas \ram_rom_data_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[8]~8_combout ),
	.asdata(ram_rom_data_reg_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N29
dffeas \ram_rom_data_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[9]~9_combout ),
	.asdata(ram_rom_data_reg_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N19
dffeas \ram_rom_data_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[10]~10_combout ),
	.asdata(ram_rom_data_reg_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N13
dffeas \ram_rom_data_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[11]~11_combout ),
	.asdata(ram_rom_data_reg_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N27
dffeas \ram_rom_data_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[12]~12_combout ),
	.asdata(ram_rom_data_reg_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N25
dffeas \ram_rom_data_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[13]~13_combout ),
	.asdata(ram_rom_data_reg_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N25
dffeas \ram_rom_data_reg[14] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[14]~14_combout ),
	.asdata(ram_rom_data_reg_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_14),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[14] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N15
dffeas \ram_rom_data_reg[15] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[15]~15_combout ),
	.asdata(ram_rom_data_reg_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_15),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[15] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N29
dffeas \ram_rom_data_reg[16] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[16]~16_combout ),
	.asdata(ram_rom_data_reg_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_16),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[16] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N11
dffeas \ram_rom_data_reg[17] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[17]~17_combout ),
	.asdata(ram_rom_data_reg_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_17),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[17] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N9
dffeas \ram_rom_data_reg[18] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[18]~18_combout ),
	.asdata(ram_rom_data_reg_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_18),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[18] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N23
dffeas \ram_rom_data_reg[19] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[19]~19_combout ),
	.asdata(ram_rom_data_reg_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_19),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[19] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N17
dffeas \ram_rom_data_reg[20] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[20]~20_combout ),
	.asdata(ram_rom_data_reg_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_20),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[20] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N31
dffeas \ram_rom_data_reg[21] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[21]~21_combout ),
	.asdata(ram_rom_data_reg_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_21),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[21] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N13
dffeas \ram_rom_data_reg[22] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[22]~22_combout ),
	.asdata(ram_rom_data_reg_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_22),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[22] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N27
dffeas \ram_rom_data_reg[23] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[23]~23_combout ),
	.asdata(ram_rom_data_reg_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_23),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[23] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N5
dffeas \ram_rom_data_reg[24] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[24]~24_combout ),
	.asdata(ram_rom_data_reg_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_24),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[24] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N15
dffeas \ram_rom_data_reg[25] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[25]~25_combout ),
	.asdata(ram_rom_data_reg_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_25),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[25] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N29
dffeas \ram_rom_data_reg[26] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[26]~26_combout ),
	.asdata(ram_rom_data_reg_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_26),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[26] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N23
dffeas \ram_rom_data_reg[27] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[27]~27_combout ),
	.asdata(ram_rom_data_reg_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_27),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[27] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N25
dffeas \ram_rom_data_reg[28] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[28]~28_combout ),
	.asdata(ram_rom_data_reg_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_28),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[28] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N7
dffeas \ram_rom_data_reg[29] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[29]~29_combout ),
	.asdata(ram_rom_data_reg_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_29),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[29] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N17
dffeas \ram_rom_data_reg[30] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[30]~30_combout ),
	.asdata(ram_rom_data_reg_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_30),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[30] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N19
dffeas \ram_rom_data_reg[31] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[31]~31_combout ),
	.asdata(altera_internal_jtag),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[0]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_31),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[31] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y34_N23
dffeas \ir_loaded_address_reg[0] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[0] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y34_N9
dffeas \ir_loaded_address_reg[1] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[1] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y34_N19
dffeas \ir_loaded_address_reg[2] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[2] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y34_N17
dffeas \ir_loaded_address_reg[3] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[3] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N30
cycloneive_lcell_comb \tdo~1 (
	.dataa(gnd),
	.datab(\tdo~0_combout ),
	.datac(ir_in[0]),
	.datad(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.cin(gnd),
	.combout(tdo),
	.cout());
// synopsys translate_off
defparam \tdo~1 .lut_mask = 16'hFC0C;
defparam \tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N24
cycloneive_lcell_comb \sdr~0 (
	.dataa(gnd),
	.datab(node_ena_1),
	.datac(virtual_ir_scan_reg),
	.datad(gnd),
	.cin(gnd),
	.combout(sdr),
	.cout());
// synopsys translate_off
defparam \sdr~0 .lut_mask = 16'h0C0C;
defparam \sdr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N12
cycloneive_lcell_comb \is_in_use_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(is_in_use_reg1),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\is_in_use_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \is_in_use_reg~0 .lut_mask = 16'h00F0;
defparam \is_in_use_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N0
cycloneive_lcell_comb \ram_rom_data_reg[0]~0 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a32),
	.datac(gnd),
	.datad(ram_block3a0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~0 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N8
cycloneive_lcell_comb \Add1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h55AA;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N10
cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h3C3F;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N4
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[1]~5 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datab(\Equal1~1_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\Add1~2_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1]~5 .lut_mask = 16'h3A10;
defparam \ram_rom_data_shift_cntr_reg[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N5
dffeas \ram_rom_data_shift_cntr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[1]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N12
cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'hC30C;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N2
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~4 (
	.dataa(irf_reg_2_1),
	.datab(irf_reg_1_1),
	.datac(state_4),
	.datad(sdr),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~4 .lut_mask = 16'hE000;
defparam \ram_rom_data_shift_cntr_reg[5]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N20
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~11 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(\Equal1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~11 .lut_mask = 16'h007F;
defparam \ram_rom_data_shift_cntr_reg[5]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N0
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[2]~9 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~4_combout ),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2]~9 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[2]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N1
dffeas \ram_rom_data_shift_cntr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[2]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N16
cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'hC30C;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N24
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[4]~7 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~8_combout ),
	.datac(ram_rom_data_shift_cntr_reg[4]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4]~7 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N25
dffeas \ram_rom_data_shift_cntr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[4]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N18
cycloneive_lcell_comb \Add1~10 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h5A5A;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N26
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~10 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~10_combout ),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~10 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[5]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N27
dffeas \ram_rom_data_shift_cntr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[5]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N28
cycloneive_lcell_comb \Equal1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(ram_rom_data_shift_cntr_reg[2]),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0800;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N22
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[0]~6 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\Add1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0]~6 .lut_mask = 16'hF444;
defparam \ram_rom_data_shift_cntr_reg[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N23
dffeas \ram_rom_data_shift_cntr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[0]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N2
cycloneive_lcell_comb \Equal1~1 (
	.dataa(gnd),
	.datab(\Equal1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'hC0C0;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N12
cycloneive_lcell_comb \process_0~2 (
	.dataa(\Equal1~1_combout ),
	.datab(irf_reg_1_1),
	.datac(ir_in[3]),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\process_0~2_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~2 .lut_mask = 16'h070F;
defparam \process_0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N20
cycloneive_lcell_comb \ram_rom_data_reg[0]~32 (
	.dataa(\process_0~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~32_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~32 .lut_mask = 16'hFF55;
defparam \ram_rom_data_reg[0]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N4
cycloneive_lcell_comb \ram_rom_addr_reg[0]~14 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[0]~14_combout ),
	.cout(\ram_rom_addr_reg[0]~15 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[0]~14 .lut_mask = 16'h33CC;
defparam \ram_rom_addr_reg[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N6
cycloneive_lcell_comb \ram_rom_addr_reg[1]~16 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[0]~15 ),
	.combout(\ram_rom_addr_reg[1]~16_combout ),
	.cout(\ram_rom_addr_reg[1]~17 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~16 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[1]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N8
cycloneive_lcell_comb \ram_rom_addr_reg[2]~18 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[1]~17 ),
	.combout(\ram_rom_addr_reg[2]~18_combout ),
	.cout(\ram_rom_addr_reg[2]~19 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~18 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[2]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N10
cycloneive_lcell_comb \ram_rom_addr_reg[3]~20 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[2]~19 ),
	.combout(\ram_rom_addr_reg[3]~20_combout ),
	.cout(\ram_rom_addr_reg[3]~21 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[3]~20 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[3]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N12
cycloneive_lcell_comb \ram_rom_addr_reg[4]~22 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[3]~21 ),
	.combout(\ram_rom_addr_reg[4]~22_combout ),
	.cout(\ram_rom_addr_reg[4]~23 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~22 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[4]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N14
cycloneive_lcell_comb \ram_rom_addr_reg[5]~24 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[4]~23 ),
	.combout(\ram_rom_addr_reg[5]~24_combout ),
	.cout(\ram_rom_addr_reg[5]~25 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~24 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[5]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N16
cycloneive_lcell_comb \ram_rom_addr_reg[6]~26 (
	.dataa(ram_rom_addr_reg_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[5]~25 ),
	.combout(\ram_rom_addr_reg[6]~26_combout ),
	.cout(\ram_rom_addr_reg[6]~27 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~26 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[6]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N18
cycloneive_lcell_comb \ram_rom_addr_reg[7]~28 (
	.dataa(ram_rom_addr_reg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[6]~27 ),
	.combout(\ram_rom_addr_reg[7]~28_combout ),
	.cout(\ram_rom_addr_reg[7]~29 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~28 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[7]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N20
cycloneive_lcell_comb \ram_rom_addr_reg[8]~30 (
	.dataa(ram_rom_addr_reg_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[7]~29 ),
	.combout(\ram_rom_addr_reg[8]~30_combout ),
	.cout(\ram_rom_addr_reg[8]~31 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[8]~30 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[8]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N22
cycloneive_lcell_comb \ram_rom_addr_reg[9]~32 (
	.dataa(ram_rom_addr_reg_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[8]~31 ),
	.combout(\ram_rom_addr_reg[9]~32_combout ),
	.cout(\ram_rom_addr_reg[9]~33 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~32 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[9]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N24
cycloneive_lcell_comb \ram_rom_addr_reg[10]~34 (
	.dataa(ram_rom_addr_reg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[9]~33 ),
	.combout(\ram_rom_addr_reg[10]~34_combout ),
	.cout(\ram_rom_addr_reg[10]~35 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[10]~34 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[10]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N26
cycloneive_lcell_comb \ram_rom_addr_reg[11]~36 (
	.dataa(ram_rom_addr_reg_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[10]~35 ),
	.combout(\ram_rom_addr_reg[11]~36_combout ),
	.cout(\ram_rom_addr_reg[11]~37 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[11]~36 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[11]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N28
cycloneive_lcell_comb \ram_rom_addr_reg[12]~38 (
	.dataa(ram_rom_addr_reg_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[11]~37 ),
	.combout(\ram_rom_addr_reg[12]~38_combout ),
	.cout(\ram_rom_addr_reg[12]~39 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[12]~38 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[12]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N30
cycloneive_lcell_comb \ram_rom_addr_reg[13]~40 (
	.dataa(ram_rom_addr_reg_13),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\ram_rom_addr_reg[12]~39 ),
	.combout(\ram_rom_addr_reg[13]~40_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[13]~40 .lut_mask = 16'h5A5A;
defparam \ram_rom_addr_reg[13]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N2
cycloneive_lcell_comb \process_0~3 (
	.dataa(state_4),
	.datab(virtual_ir_scan_reg),
	.datac(node_ena_1),
	.datad(ir_in[3]),
	.cin(gnd),
	.combout(\process_0~3_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~3 .lut_mask = 16'h2000;
defparam \process_0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N26
cycloneive_lcell_comb \ram_rom_addr_reg[9]~42 (
	.dataa(\Equal1~1_combout ),
	.datab(irf_reg_1_1),
	.datac(\process_0~3_combout ),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[9]~42_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~42 .lut_mask = 16'hF0F8;
defparam \ram_rom_addr_reg[9]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N8
cycloneive_lcell_comb \ram_rom_addr_reg[9]~43 (
	.dataa(state_8),
	.datab(sdr),
	.datac(\ram_rom_addr_reg[9]~42_combout ),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[9]~43_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~43 .lut_mask = 16'hF8F0;
defparam \ram_rom_addr_reg[9]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N16
cycloneive_lcell_comb \ram_rom_data_reg[1]~1 (
	.dataa(ram_block3a1),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a33),
	.cin(gnd),
	.combout(\ram_rom_data_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[1]~1 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N22
cycloneive_lcell_comb \ram_rom_data_reg[2]~2 (
	.dataa(ram_block3a2),
	.datab(ram_block3a34),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[2]~2 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N8
cycloneive_lcell_comb \ram_rom_data_reg[3]~3 (
	.dataa(ram_block3a35),
	.datab(ram_block3a3),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[3]~3 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N26
cycloneive_lcell_comb \ram_rom_data_reg[4]~4 (
	.dataa(ram_block3a4),
	.datab(ram_block3a36),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[4]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[4]~4 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N24
cycloneive_lcell_comb \ram_rom_data_reg[5]~5 (
	.dataa(ram_block3a5),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a37),
	.cin(gnd),
	.combout(\ram_rom_data_reg[5]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[5]~5 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N14
cycloneive_lcell_comb \ram_rom_data_reg[6]~6 (
	.dataa(ram_block3a38),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a6),
	.cin(gnd),
	.combout(\ram_rom_data_reg[6]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[6]~6 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N20
cycloneive_lcell_comb \ram_rom_data_reg[7]~7 (
	.dataa(ram_block3a7),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a39),
	.cin(gnd),
	.combout(\ram_rom_data_reg[7]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[7]~7 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N30
cycloneive_lcell_comb \ram_rom_data_reg[8]~8 (
	.dataa(ram_block3a8),
	.datab(ram_block3a40),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[8]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[8]~8 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N28
cycloneive_lcell_comb \ram_rom_data_reg[9]~9 (
	.dataa(ram_block3a41),
	.datab(ram_block3a9),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[9]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[9]~9 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N18
cycloneive_lcell_comb \ram_rom_data_reg[10]~10 (
	.dataa(ram_block3a10),
	.datab(ram_block3a42),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[10]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[10]~10 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N12
cycloneive_lcell_comb \ram_rom_data_reg[11]~11 (
	.dataa(ram_block3a11),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a43),
	.cin(gnd),
	.combout(\ram_rom_data_reg[11]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[11]~11 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N26
cycloneive_lcell_comb \ram_rom_data_reg[12]~12 (
	.dataa(ram_block3a12),
	.datab(ram_block3a44),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~12 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N24
cycloneive_lcell_comb \ram_rom_data_reg[13]~13 (
	.dataa(ram_block3a13),
	.datab(ram_block3a45),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[13]~13_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[13]~13 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N24
cycloneive_lcell_comb \ram_rom_data_reg[14]~14 (
	.dataa(ram_block3a14),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a46),
	.cin(gnd),
	.combout(\ram_rom_data_reg[14]~14_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[14]~14 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N14
cycloneive_lcell_comb \ram_rom_data_reg[15]~15 (
	.dataa(ram_block3a15),
	.datab(ram_block3a47),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[15]~15_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[15]~15 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N28
cycloneive_lcell_comb \ram_rom_data_reg[16]~16 (
	.dataa(ram_block3a16),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a48),
	.cin(gnd),
	.combout(\ram_rom_data_reg[16]~16_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[16]~16 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N10
cycloneive_lcell_comb \ram_rom_data_reg[17]~17 (
	.dataa(ram_block3a17),
	.datab(ram_block3a49),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[17]~17_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[17]~17 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N8
cycloneive_lcell_comb \ram_rom_data_reg[18]~18 (
	.dataa(ram_block3a18),
	.datab(ram_block3a50),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[18]~18_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[18]~18 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N22
cycloneive_lcell_comb \ram_rom_data_reg[19]~19 (
	.dataa(ram_block3a19),
	.datab(ram_block3a51),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[19]~19_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[19]~19 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N16
cycloneive_lcell_comb \ram_rom_data_reg[20]~20 (
	.dataa(ram_block3a52),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a20),
	.cin(gnd),
	.combout(\ram_rom_data_reg[20]~20_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[20]~20 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N30
cycloneive_lcell_comb \ram_rom_data_reg[21]~21 (
	.dataa(ram_block3a53),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a21),
	.cin(gnd),
	.combout(\ram_rom_data_reg[21]~21_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[21]~21 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N12
cycloneive_lcell_comb \ram_rom_data_reg[22]~22 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a54),
	.datac(gnd),
	.datad(ram_block3a22),
	.cin(gnd),
	.combout(\ram_rom_data_reg[22]~22_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[22]~22 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N26
cycloneive_lcell_comb \ram_rom_data_reg[23]~23 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a23),
	.datac(gnd),
	.datad(ram_block3a55),
	.cin(gnd),
	.combout(\ram_rom_data_reg[23]~23_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[23]~23 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N4
cycloneive_lcell_comb \ram_rom_data_reg[24]~24 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a56),
	.datac(gnd),
	.datad(ram_block3a24),
	.cin(gnd),
	.combout(\ram_rom_data_reg[24]~24_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[24]~24 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N14
cycloneive_lcell_comb \ram_rom_data_reg[25]~25 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a57),
	.datac(gnd),
	.datad(ram_block3a25),
	.cin(gnd),
	.combout(\ram_rom_data_reg[25]~25_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[25]~25 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N28
cycloneive_lcell_comb \ram_rom_data_reg[26]~26 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a26),
	.datac(gnd),
	.datad(ram_block3a58),
	.cin(gnd),
	.combout(\ram_rom_data_reg[26]~26_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[26]~26 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N22
cycloneive_lcell_comb \ram_rom_data_reg[27]~27 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a59),
	.datac(gnd),
	.datad(ram_block3a27),
	.cin(gnd),
	.combout(\ram_rom_data_reg[27]~27_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[27]~27 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N24
cycloneive_lcell_comb \ram_rom_data_reg[28]~28 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a28),
	.datac(gnd),
	.datad(ram_block3a60),
	.cin(gnd),
	.combout(\ram_rom_data_reg[28]~28_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[28]~28 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N6
cycloneive_lcell_comb \ram_rom_data_reg[29]~29 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a29),
	.datac(gnd),
	.datad(ram_block3a61),
	.cin(gnd),
	.combout(\ram_rom_data_reg[29]~29_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[29]~29 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N16
cycloneive_lcell_comb \ram_rom_data_reg[30]~30 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a30),
	.datac(gnd),
	.datad(ram_block3a62),
	.cin(gnd),
	.combout(\ram_rom_data_reg[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[30]~30 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N18
cycloneive_lcell_comb \ram_rom_data_reg[31]~31 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a31),
	.datac(gnd),
	.datad(ram_block3a63),
	.cin(gnd),
	.combout(\ram_rom_data_reg[31]~31_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[31]~31 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N22
cycloneive_lcell_comb \ir_loaded_address_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(ram_rom_addr_reg_0),
	.datad(gnd),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[0]~feeder .lut_mask = 16'hF0F0;
defparam \ir_loaded_address_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N30
cycloneive_lcell_comb \process_0~0 (
	.dataa(gnd),
	.datab(irf_reg_4_1),
	.datac(ir_in[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\process_0~0_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~0 .lut_mask = 16'hFCFC;
defparam \process_0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N0
cycloneive_lcell_comb \process_0~1 (
	.dataa(virtual_ir_scan_reg),
	.datab(node_ena_1),
	.datac(state_5),
	.datad(ir_in[3]),
	.cin(gnd),
	.combout(\process_0~1_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~1 .lut_mask = 16'h4000;
defparam \process_0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N8
cycloneive_lcell_comb \ir_loaded_address_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_1),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N18
cycloneive_lcell_comb \ir_loaded_address_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_2),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N16
cycloneive_lcell_comb \ir_loaded_address_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_3),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N14
cycloneive_lcell_comb \bypass_reg_out~0 (
	.dataa(gnd),
	.datab(node_ena_1),
	.datac(\bypass_reg_out~q ),
	.datad(altera_internal_jtag),
	.cin(gnd),
	.combout(\bypass_reg_out~0_combout ),
	.cout());
// synopsys translate_off
defparam \bypass_reg_out~0 .lut_mask = 16'hFC30;
defparam \bypass_reg_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N15
dffeas bypass_reg_out(
	.clk(raw_tck),
	.d(\bypass_reg_out~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bypass_reg_out~q ),
	.prn(vcc));
// synopsys translate_off
defparam bypass_reg_out.is_wysiwyg = "true";
defparam bypass_reg_out.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N28
cycloneive_lcell_comb \tdo~0 (
	.dataa(\bypass_reg_out~q ),
	.datab(irf_reg_1_1),
	.datac(ram_rom_data_reg_0),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \tdo~0 .lut_mask = 16'hF0E2;
defparam \tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_rom_sr (
	WORD_SR_0,
	sdr,
	altera_internal_jtag,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	TCK,
	devpor,
	devclrn,
	devoe);
output 	WORD_SR_0;
input 	sdr;
input 	altera_internal_jtag;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	TCK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \word_counter[3]~15_combout ;
wire \WORD_SR~3_combout ;
wire \WORD_SR~7_combout ;
wire \WORD_SR~8_combout ;
wire \WORD_SR~13_combout ;
wire \WORD_SR~14_combout ;
wire \WORD_SR~15_combout ;
wire \word_counter[0]~7_combout ;
wire \word_counter[0]~8 ;
wire \word_counter[1]~10 ;
wire \word_counter[2]~11_combout ;
wire \clear_signal~combout ;
wire \word_counter[0]~14_combout ;
wire \word_counter[2]~12 ;
wire \word_counter[3]~16 ;
wire \word_counter[4]~17_combout ;
wire \word_counter[1]~9_combout ;
wire \word_counter[0]~13_combout ;
wire \word_counter[0]~19_combout ;
wire \WORD_SR~2_combout ;
wire \WORD_SR~4_combout ;
wire \WORD_SR~10_combout ;
wire \WORD_SR~11_combout ;
wire \WORD_SR~12_combout ;
wire \WORD_SR[1]~6_combout ;
wire \WORD_SR~9_combout ;
wire \WORD_SR~5_combout ;
wire [4:0] word_counter;
wire [3:0] WORD_SR;


// Location: FF_X41_Y34_N11
dffeas \word_counter[3] (
	.clk(TCK),
	.d(\word_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[3]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[3] .is_wysiwyg = "true";
defparam \word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N10
cycloneive_lcell_comb \word_counter[3]~15 (
	.dataa(word_counter[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[2]~12 ),
	.combout(\word_counter[3]~15_combout ),
	.cout(\word_counter[3]~16 ));
// synopsys translate_off
defparam \word_counter[3]~15 .lut_mask = 16'h5A5F;
defparam \word_counter[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N22
cycloneive_lcell_comb \WORD_SR~3 (
	.dataa(word_counter[4]),
	.datab(word_counter[0]),
	.datac(word_counter[2]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~3_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~3 .lut_mask = 16'hBA02;
defparam \WORD_SR~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N0
cycloneive_lcell_comb \WORD_SR~7 (
	.dataa(state_4),
	.datab(word_counter[0]),
	.datac(word_counter[1]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~7 .lut_mask = 16'h1011;
defparam \WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N10
cycloneive_lcell_comb \WORD_SR~8 (
	.dataa(word_counter[3]),
	.datab(\WORD_SR~7_combout ),
	.datac(gnd),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~8 .lut_mask = 16'h0044;
defparam \WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N27
dffeas \WORD_SR[3] (
	.clk(TCK),
	.d(\WORD_SR~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[1]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[3]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[3] .is_wysiwyg = "true";
defparam \WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N24
cycloneive_lcell_comb \WORD_SR~13 (
	.dataa(word_counter[3]),
	.datab(word_counter[4]),
	.datac(word_counter[2]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~13 .lut_mask = 16'h2000;
defparam \WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N20
cycloneive_lcell_comb \WORD_SR~14 (
	.dataa(state_4),
	.datab(altera_internal_jtag),
	.datac(word_counter[0]),
	.datad(\WORD_SR~13_combout ),
	.cin(gnd),
	.combout(\WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~14 .lut_mask = 16'h8D88;
defparam \WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N26
cycloneive_lcell_comb \WORD_SR~15 (
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(state_8),
	.datad(\WORD_SR~14_combout ),
	.cin(gnd),
	.combout(\WORD_SR~15_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~15 .lut_mask = 16'h5F00;
defparam \WORD_SR~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N25
dffeas \WORD_SR[0] (
	.clk(TCK),
	.d(\WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[1]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR_0),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[0] .is_wysiwyg = "true";
defparam \WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N4
cycloneive_lcell_comb \word_counter[0]~7 (
	.dataa(gnd),
	.datab(word_counter[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\word_counter[0]~7_combout ),
	.cout(\word_counter[0]~8 ));
// synopsys translate_off
defparam \word_counter[0]~7 .lut_mask = 16'h33CC;
defparam \word_counter[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N6
cycloneive_lcell_comb \word_counter[1]~9 (
	.dataa(word_counter[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[0]~8 ),
	.combout(\word_counter[1]~9_combout ),
	.cout(\word_counter[1]~10 ));
// synopsys translate_off
defparam \word_counter[1]~9 .lut_mask = 16'h5A5F;
defparam \word_counter[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N8
cycloneive_lcell_comb \word_counter[2]~11 (
	.dataa(gnd),
	.datab(word_counter[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[1]~10 ),
	.combout(\word_counter[2]~11_combout ),
	.cout(\word_counter[2]~12 ));
// synopsys translate_off
defparam \word_counter[2]~11 .lut_mask = 16'hC30C;
defparam \word_counter[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N16
cycloneive_lcell_comb clear_signal(
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(state_8),
	.datad(gnd),
	.cin(gnd),
	.combout(\clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam clear_signal.lut_mask = 16'hA0A0;
defparam clear_signal.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N12
cycloneive_lcell_comb \word_counter[0]~14 (
	.dataa(sdr),
	.datab(state_3),
	.datac(state_4),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\word_counter[0]~14_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[0]~14 .lut_mask = 16'hFF08;
defparam \word_counter[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y34_N9
dffeas \word_counter[2] (
	.clk(TCK),
	.d(\word_counter[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[2]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[2] .is_wysiwyg = "true";
defparam \word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N12
cycloneive_lcell_comb \word_counter[4]~17 (
	.dataa(word_counter[4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\word_counter[3]~16 ),
	.combout(\word_counter[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~17 .lut_mask = 16'hA5A5;
defparam \word_counter[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X41_Y34_N13
dffeas \word_counter[4] (
	.clk(TCK),
	.d(\word_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[4]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[4] .is_wysiwyg = "true";
defparam \word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N7
dffeas \word_counter[1] (
	.clk(TCK),
	.d(\word_counter[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[1]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[1] .is_wysiwyg = "true";
defparam \word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N18
cycloneive_lcell_comb \word_counter[0]~13 (
	.dataa(word_counter[3]),
	.datab(word_counter[4]),
	.datac(word_counter[1]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\word_counter[0]~13_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[0]~13 .lut_mask = 16'hFBFF;
defparam \word_counter[0]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N6
cycloneive_lcell_comb \word_counter[0]~19 (
	.dataa(virtual_ir_scan_reg),
	.datab(state_8),
	.datac(word_counter[0]),
	.datad(\word_counter[0]~13_combout ),
	.cin(gnd),
	.combout(\word_counter[0]~19_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[0]~19 .lut_mask = 16'h888F;
defparam \word_counter[0]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y34_N5
dffeas \word_counter[0] (
	.clk(TCK),
	.d(\word_counter[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[0]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[0] .is_wysiwyg = "true";
defparam \word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N0
cycloneive_lcell_comb \WORD_SR~2 (
	.dataa(word_counter[3]),
	.datab(word_counter[4]),
	.datac(word_counter[2]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~2_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~2 .lut_mask = 16'h2025;
defparam \WORD_SR~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N14
cycloneive_lcell_comb \WORD_SR~4 (
	.dataa(\WORD_SR~3_combout ),
	.datab(gnd),
	.datac(word_counter[0]),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~4_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~4 .lut_mask = 16'hAAA0;
defparam \WORD_SR~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N28
cycloneive_lcell_comb \WORD_SR~10 (
	.dataa(word_counter[4]),
	.datab(word_counter[0]),
	.datac(word_counter[2]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~10 .lut_mask = 16'hCABA;
defparam \WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N2
cycloneive_lcell_comb \WORD_SR~11 (
	.dataa(gnd),
	.datab(\WORD_SR~10_combout ),
	.datac(word_counter[0]),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~11 .lut_mask = 16'hC3C0;
defparam \WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N28
cycloneive_lcell_comb \WORD_SR~12 (
	.dataa(WORD_SR[3]),
	.datab(\clear_signal~combout ),
	.datac(state_4),
	.datad(\WORD_SR~11_combout ),
	.cin(gnd),
	.combout(\WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~12 .lut_mask = 16'h2320;
defparam \WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N22
cycloneive_lcell_comb \WORD_SR[1]~6 (
	.dataa(sdr),
	.datab(state_3),
	.datac(state_4),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR[1]~6_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR[1]~6 .lut_mask = 16'hFFA8;
defparam \WORD_SR[1]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N29
dffeas \WORD_SR[2] (
	.clk(TCK),
	.d(\WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[1]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[2]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[2] .is_wysiwyg = "true";
defparam \WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N2
cycloneive_lcell_comb \WORD_SR~9 (
	.dataa(\WORD_SR~8_combout ),
	.datab(WORD_SR[2]),
	.datac(state_4),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~9 .lut_mask = 16'h00EA;
defparam \WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N3
dffeas \WORD_SR[1] (
	.clk(TCK),
	.d(\WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[1]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[1]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[1] .is_wysiwyg = "true";
defparam \WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N24
cycloneive_lcell_comb \WORD_SR~5 (
	.dataa(\WORD_SR~4_combout ),
	.datab(WORD_SR[1]),
	.datac(state_4),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR~5_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~5 .lut_mask = 16'h00CA;
defparam \WORD_SR~5 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule
